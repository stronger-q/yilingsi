module ORB_BRIEF(
    input                               i_clk,

    interface_windows.i_window     i_window,

    output    [255:0]                   o_brief
    );

logic [7:0] PA_000;
logic [7:0] PB_000;
logic [7:0] PA_001;
logic [7:0] PB_001;
logic [7:0] PA_002;
logic [7:0] PB_002;
logic [7:0] PA_003;
logic [7:0] PB_003;
logic [7:0] PA_004;
logic [7:0] PB_004;
logic [7:0] PA_005;
logic [7:0] PB_005;
logic [7:0] PA_006;
logic [7:0] PB_006;
logic [7:0] PA_007;
logic [7:0] PB_007;
logic [7:0] PA_008;
logic [7:0] PB_008;
logic [7:0] PA_009;
logic [7:0] PB_009;
logic [7:0] PA_010;
logic [7:0] PB_010;
logic [7:0] PA_011;
logic [7:0] PB_011;
logic [7:0] PA_012;
logic [7:0] PB_012;
logic [7:0] PA_013;
logic [7:0] PB_013;
logic [7:0] PA_014;
logic [7:0] PB_014;
logic [7:0] PA_015;
logic [7:0] PB_015;
logic [7:0] PA_016;
logic [7:0] PB_016;
logic [7:0] PA_017;
logic [7:0] PB_017;
logic [7:0] PA_018;
logic [7:0] PB_018;
logic [7:0] PA_019;
logic [7:0] PB_019;
logic [7:0] PA_020;
logic [7:0] PB_020;
logic [7:0] PA_021;
logic [7:0] PB_021;
logic [7:0] PA_022;
logic [7:0] PB_022;
logic [7:0] PA_023;
logic [7:0] PB_023;
logic [7:0] PA_024;
logic [7:0] PB_024;
logic [7:0] PA_025;
logic [7:0] PB_025;
logic [7:0] PA_026;
logic [7:0] PB_026;
logic [7:0] PA_027;
logic [7:0] PB_027;
logic [7:0] PA_028;
logic [7:0] PB_028;
logic [7:0] PA_029;
logic [7:0] PB_029;
logic [7:0] PA_030;
logic [7:0] PB_030;
logic [7:0] PA_031;
logic [7:0] PB_031;
logic [7:0] PA_032;
logic [7:0] PB_032;
logic [7:0] PA_033;
logic [7:0] PB_033;
logic [7:0] PA_034;
logic [7:0] PB_034;
logic [7:0] PA_035;
logic [7:0] PB_035;
logic [7:0] PA_036;
logic [7:0] PB_036;
logic [7:0] PA_037;
logic [7:0] PB_037;
logic [7:0] PA_038;
logic [7:0] PB_038;
logic [7:0] PA_039;
logic [7:0] PB_039;
logic [7:0] PA_040;
logic [7:0] PB_040;
logic [7:0] PA_041;
logic [7:0] PB_041;
logic [7:0] PA_042;
logic [7:0] PB_042;
logic [7:0] PA_043;
logic [7:0] PB_043;
logic [7:0] PA_044;
logic [7:0] PB_044;
logic [7:0] PA_045;
logic [7:0] PB_045;
logic [7:0] PA_046;
logic [7:0] PB_046;
logic [7:0] PA_047;
logic [7:0] PB_047;
logic [7:0] PA_048;
logic [7:0] PB_048;
logic [7:0] PA_049;
logic [7:0] PB_049;
logic [7:0] PA_050;
logic [7:0] PB_050;
logic [7:0] PA_051;
logic [7:0] PB_051;
logic [7:0] PA_052;
logic [7:0] PB_052;
logic [7:0] PA_053;
logic [7:0] PB_053;
logic [7:0] PA_054;
logic [7:0] PB_054;
logic [7:0] PA_055;
logic [7:0] PB_055;
logic [7:0] PA_056;
logic [7:0] PB_056;
logic [7:0] PA_057;
logic [7:0] PB_057;
logic [7:0] PA_058;
logic [7:0] PB_058;
logic [7:0] PA_059;
logic [7:0] PB_059;
logic [7:0] PA_060;
logic [7:0] PB_060;
logic [7:0] PA_061;
logic [7:0] PB_061;
logic [7:0] PA_062;
logic [7:0] PB_062;
logic [7:0] PA_063;
logic [7:0] PB_063;
logic [7:0] PA_064;
logic [7:0] PB_064;
logic [7:0] PA_065;
logic [7:0] PB_065;
logic [7:0] PA_066;
logic [7:0] PB_066;
logic [7:0] PA_067;
logic [7:0] PB_067;
logic [7:0] PA_068;
logic [7:0] PB_068;
logic [7:0] PA_069;
logic [7:0] PB_069;
logic [7:0] PA_070;
logic [7:0] PB_070;
logic [7:0] PA_071;
logic [7:0] PB_071;
logic [7:0] PA_072;
logic [7:0] PB_072;
logic [7:0] PA_073;
logic [7:0] PB_073;
logic [7:0] PA_074;
logic [7:0] PB_074;
logic [7:0] PA_075;
logic [7:0] PB_075;
logic [7:0] PA_076;
logic [7:0] PB_076;
logic [7:0] PA_077;
logic [7:0] PB_077;
logic [7:0] PA_078;
logic [7:0] PB_078;
logic [7:0] PA_079;
logic [7:0] PB_079;
logic [7:0] PA_080;
logic [7:0] PB_080;
logic [7:0] PA_081;
logic [7:0] PB_081;
logic [7:0] PA_082;
logic [7:0] PB_082;
logic [7:0] PA_083;
logic [7:0] PB_083;
logic [7:0] PA_084;
logic [7:0] PB_084;
logic [7:0] PA_085;
logic [7:0] PB_085;
logic [7:0] PA_086;
logic [7:0] PB_086;
logic [7:0] PA_087;
logic [7:0] PB_087;
logic [7:0] PA_088;
logic [7:0] PB_088;
logic [7:0] PA_089;
logic [7:0] PB_089;
logic [7:0] PA_090;
logic [7:0] PB_090;
logic [7:0] PA_091;
logic [7:0] PB_091;
logic [7:0] PA_092;
logic [7:0] PB_092;
logic [7:0] PA_093;
logic [7:0] PB_093;
logic [7:0] PA_094;
logic [7:0] PB_094;
logic [7:0] PA_095;
logic [7:0] PB_095;
logic [7:0] PA_096;
logic [7:0] PB_096;
logic [7:0] PA_097;
logic [7:0] PB_097;
logic [7:0] PA_098;
logic [7:0] PB_098;
logic [7:0] PA_099;
logic [7:0] PB_099;
logic [7:0] PA_100;
logic [7:0] PB_100;
logic [7:0] PA_101;
logic [7:0] PB_101;
logic [7:0] PA_102;
logic [7:0] PB_102;
logic [7:0] PA_103;
logic [7:0] PB_103;
logic [7:0] PA_104;
logic [7:0] PB_104;
logic [7:0] PA_105;
logic [7:0] PB_105;
logic [7:0] PA_106;
logic [7:0] PB_106;
logic [7:0] PA_107;
logic [7:0] PB_107;
logic [7:0] PA_108;
logic [7:0] PB_108;
logic [7:0] PA_109;
logic [7:0] PB_109;
logic [7:0] PA_110;
logic [7:0] PB_110;
logic [7:0] PA_111;
logic [7:0] PB_111;
logic [7:0] PA_112;
logic [7:0] PB_112;
logic [7:0] PA_113;
logic [7:0] PB_113;
logic [7:0] PA_114;
logic [7:0] PB_114;
logic [7:0] PA_115;
logic [7:0] PB_115;
logic [7:0] PA_116;
logic [7:0] PB_116;
logic [7:0] PA_117;
logic [7:0] PB_117;
logic [7:0] PA_118;
logic [7:0] PB_118;
logic [7:0] PA_119;
logic [7:0] PB_119;
logic [7:0] PA_120;
logic [7:0] PB_120;
logic [7:0] PA_121;
logic [7:0] PB_121;
logic [7:0] PA_122;
logic [7:0] PB_122;
logic [7:0] PA_123;
logic [7:0] PB_123;
logic [7:0] PA_124;
logic [7:0] PB_124;
logic [7:0] PA_125;
logic [7:0] PB_125;
logic [7:0] PA_126;
logic [7:0] PB_126;
logic [7:0] PA_127;
logic [7:0] PB_127;
logic [7:0] PA_128;
logic [7:0] PB_128;
logic [7:0] PA_129;
logic [7:0] PB_129;
logic [7:0] PA_130;
logic [7:0] PB_130;
logic [7:0] PA_131;
logic [7:0] PB_131;
logic [7:0] PA_132;
logic [7:0] PB_132;
logic [7:0] PA_133;
logic [7:0] PB_133;
logic [7:0] PA_134;
logic [7:0] PB_134;
logic [7:0] PA_135;
logic [7:0] PB_135;
logic [7:0] PA_136;
logic [7:0] PB_136;
logic [7:0] PA_137;
logic [7:0] PB_137;
logic [7:0] PA_138;
logic [7:0] PB_138;
logic [7:0] PA_139;
logic [7:0] PB_139;
logic [7:0] PA_140;
logic [7:0] PB_140;
logic [7:0] PA_141;
logic [7:0] PB_141;
logic [7:0] PA_142;
logic [7:0] PB_142;
logic [7:0] PA_143;
logic [7:0] PB_143;
logic [7:0] PA_144;
logic [7:0] PB_144;
logic [7:0] PA_145;
logic [7:0] PB_145;
logic [7:0] PA_146;
logic [7:0] PB_146;
logic [7:0] PA_147;
logic [7:0] PB_147;
logic [7:0] PA_148;
logic [7:0] PB_148;
logic [7:0] PA_149;
logic [7:0] PB_149;
logic [7:0] PA_150;
logic [7:0] PB_150;
logic [7:0] PA_151;
logic [7:0] PB_151;
logic [7:0] PA_152;
logic [7:0] PB_152;
logic [7:0] PA_153;
logic [7:0] PB_153;
logic [7:0] PA_154;
logic [7:0] PB_154;
logic [7:0] PA_155;
logic [7:0] PB_155;
logic [7:0] PA_156;
logic [7:0] PB_156;
logic [7:0] PA_157;
logic [7:0] PB_157;
logic [7:0] PA_158;
logic [7:0] PB_158;
logic [7:0] PA_159;
logic [7:0] PB_159;
logic [7:0] PA_160;
logic [7:0] PB_160;
logic [7:0] PA_161;
logic [7:0] PB_161;
logic [7:0] PA_162;
logic [7:0] PB_162;
logic [7:0] PA_163;
logic [7:0] PB_163;
logic [7:0] PA_164;
logic [7:0] PB_164;
logic [7:0] PA_165;
logic [7:0] PB_165;
logic [7:0] PA_166;
logic [7:0] PB_166;
logic [7:0] PA_167;
logic [7:0] PB_167;
logic [7:0] PA_168;
logic [7:0] PB_168;
logic [7:0] PA_169;
logic [7:0] PB_169;
logic [7:0] PA_170;
logic [7:0] PB_170;
logic [7:0] PA_171;
logic [7:0] PB_171;
logic [7:0] PA_172;
logic [7:0] PB_172;
logic [7:0] PA_173;
logic [7:0] PB_173;
logic [7:0] PA_174;
logic [7:0] PB_174;
logic [7:0] PA_175;
logic [7:0] PB_175;
logic [7:0] PA_176;
logic [7:0] PB_176;
logic [7:0] PA_177;
logic [7:0] PB_177;
logic [7:0] PA_178;
logic [7:0] PB_178;
logic [7:0] PA_179;
logic [7:0] PB_179;
logic [7:0] PA_180;
logic [7:0] PB_180;
logic [7:0] PA_181;
logic [7:0] PB_181;
logic [7:0] PA_182;
logic [7:0] PB_182;
logic [7:0] PA_183;
logic [7:0] PB_183;
logic [7:0] PA_184;
logic [7:0] PB_184;
logic [7:0] PA_185;
logic [7:0] PB_185;
logic [7:0] PA_186;
logic [7:0] PB_186;
logic [7:0] PA_187;
logic [7:0] PB_187;
logic [7:0] PA_188;
logic [7:0] PB_188;
logic [7:0] PA_189;
logic [7:0] PB_189;
logic [7:0] PA_190;
logic [7:0] PB_190;
logic [7:0] PA_191;
logic [7:0] PB_191;
logic [7:0] PA_192;
logic [7:0] PB_192;
logic [7:0] PA_193;
logic [7:0] PB_193;
logic [7:0] PA_194;
logic [7:0] PB_194;
logic [7:0] PA_195;
logic [7:0] PB_195;
logic [7:0] PA_196;
logic [7:0] PB_196;
logic [7:0] PA_197;
logic [7:0] PB_197;
logic [7:0] PA_198;
logic [7:0] PB_198;
logic [7:0] PA_199;
logic [7:0] PB_199;
logic [7:0] PA_200;
logic [7:0] PB_200;
logic [7:0] PA_201;
logic [7:0] PB_201;
logic [7:0] PA_202;
logic [7:0] PB_202;
logic [7:0] PA_203;
logic [7:0] PB_203;
logic [7:0] PA_204;
logic [7:0] PB_204;
logic [7:0] PA_205;
logic [7:0] PB_205;
logic [7:0] PA_206;
logic [7:0] PB_206;
logic [7:0] PA_207;
logic [7:0] PB_207;
logic [7:0] PA_208;
logic [7:0] PB_208;
logic [7:0] PA_209;
logic [7:0] PB_209;
logic [7:0] PA_210;
logic [7:0] PB_210;
logic [7:0] PA_211;
logic [7:0] PB_211;
logic [7:0] PA_212;
logic [7:0] PB_212;
logic [7:0] PA_213;
logic [7:0] PB_213;
logic [7:0] PA_214;
logic [7:0] PB_214;
logic [7:0] PA_215;
logic [7:0] PB_215;
logic [7:0] PA_216;
logic [7:0] PB_216;
logic [7:0] PA_217;
logic [7:0] PB_217;
logic [7:0] PA_218;
logic [7:0] PB_218;
logic [7:0] PA_219;
logic [7:0] PB_219;
logic [7:0] PA_220;
logic [7:0] PB_220;
logic [7:0] PA_221;
logic [7:0] PB_221;
logic [7:0] PA_222;
logic [7:0] PB_222;
logic [7:0] PA_223;
logic [7:0] PB_223;
logic [7:0] PA_224;
logic [7:0] PB_224;
logic [7:0] PA_225;
logic [7:0] PB_225;
logic [7:0] PA_226;
logic [7:0] PB_226;
logic [7:0] PA_227;
logic [7:0] PB_227;
logic [7:0] PA_228;
logic [7:0] PB_228;
logic [7:0] PA_229;
logic [7:0] PB_229;
logic [7:0] PA_230;
logic [7:0] PB_230;
logic [7:0] PA_231;
logic [7:0] PB_231;
logic [7:0] PA_232;
logic [7:0] PB_232;
logic [7:0] PA_233;
logic [7:0] PB_233;
logic [7:0] PA_234;
logic [7:0] PB_234;
logic [7:0] PA_235;
logic [7:0] PB_235;
logic [7:0] PA_236;
logic [7:0] PB_236;
logic [7:0] PA_237;
logic [7:0] PB_237;
logic [7:0] PA_238;
logic [7:0] PB_238;
logic [7:0] PA_239;
logic [7:0] PB_239;
logic [7:0] PA_240;
logic [7:0] PB_240;
logic [7:0] PA_241;
logic [7:0] PB_241;
logic [7:0] PA_242;
logic [7:0] PB_242;
logic [7:0] PA_243;
logic [7:0] PB_243;
logic [7:0] PA_244;
logic [7:0] PB_244;
logic [7:0] PA_245;
logic [7:0] PB_245;
logic [7:0] PA_246;
logic [7:0] PB_246;
logic [7:0] PA_247;
logic [7:0] PB_247;
logic [7:0] PA_248;
logic [7:0] PB_248;
logic [7:0] PA_249;
logic [7:0] PB_249;
logic [7:0] PA_250;
logic [7:0] PB_250;
logic [7:0] PA_251;
logic [7:0] PB_251;
logic [7:0] PA_252;
logic [7:0] PB_252;
logic [7:0] PA_253;
logic [7:0] PB_253;
logic [7:0] PA_254;
logic [7:0] PB_254;
logic [7:0] PA_255;
logic [7:0] PB_255;


assign PA_000= i_window.window_12[23];
assign PB_000= i_window.window_20[24];
assign PA_001= i_window.window_17[19];
assign PB_001= i_window.window_03[22];
assign PA_002= i_window.window_24[04];
assign PB_002= i_window.window_17[07];
assign PA_003= i_window.window_03[22];
assign PB_003= i_window.window_02[27];
assign PA_004= i_window.window_02[17];
assign PB_004= i_window.window_27[17];
assign PA_005= i_window.window_08[16];
assign PB_005= i_window.window_21[16];
assign PA_006= i_window.window_05[13];
assign PB_006= i_window.window_11[13];
assign PA_007= i_window.window_02[02];
assign PB_007= i_window.window_07[04];
assign PA_008= i_window.window_12[02];
assign PB_008= i_window.window_06[03];
assign PA_009= i_window.window_19[25];
assign PB_009= i_window.window_24[26];
assign PA_010= i_window.window_07[02];
assign PB_010= i_window.window_06[07];
assign PA_011= i_window.window_22[04];
assign PB_011= i_window.window_27[06];
assign PA_012= i_window.window_22[22];
assign PB_012= i_window.window_21[27];
assign PA_013= i_window.window_10[11];
assign PB_013= i_window.window_15[12];
assign PA_014= i_window.window_17[02];
assign PB_014= i_window.window_12[03];
assign PA_015= i_window.window_15[06];
assign PB_015= i_window.window_20[08];
assign PA_016= i_window.window_09[27];
assign PB_016= i_window.window_14[27];
assign PA_017= i_window.window_21[12];
assign PB_017= i_window.window_27[13];
assign PA_018= i_window.window_02[09];
assign PB_018= i_window.window_07[11];
assign PA_019= i_window.window_02[26];
assign PB_019= i_window.window_07[27];
assign PA_020= i_window.window_22[19];
assign PB_020= i_window.window_16[20];
assign PA_021= i_window.window_12[20];
assign PB_021= i_window.window_12[25];
assign PA_022= i_window.window_08[18];
assign PB_022= i_window.window_27[21];
assign PA_023= i_window.window_08[07];
assign PB_023= i_window.window_13[09];
assign PA_024= i_window.window_26[13];
assign PB_024= i_window.window_05[14];
assign PA_025= i_window.window_27[02];
assign PB_025= i_window.window_25[07];
assign PA_026= i_window.window_18[08];
assign PB_026= i_window.window_12[10];
assign PA_027= i_window.window_17[11];
assign PB_027= i_window.window_22[12];
assign PA_028= i_window.window_03[05];
assign PB_028= i_window.window_26[09];
assign PA_029= i_window.window_03[20];
assign PB_029= i_window.window_08[21];
assign PA_030= i_window.window_09[20];
assign PB_030= i_window.window_14[22];
assign PA_031= i_window.window_15[16];
assign PB_031= i_window.window_10[19];
assign PA_032= i_window.window_26[24];
assign PB_032= i_window.window_02[26];
assign PA_033= i_window.window_22[19];
assign PB_033= i_window.window_27[19];
assign PA_034= i_window.window_14[17];
assign PB_034= i_window.window_19[19];
assign PA_035= i_window.window_03[11];
assign PB_035= i_window.window_22[13];
assign PA_036= i_window.window_10[07];
assign PB_036= i_window.window_05[08];
assign PA_037= i_window.window_26[19];
assign PB_037= i_window.window_27[24];
assign PA_038= i_window.window_07[15];
assign PB_038= i_window.window_02[16];
assign PA_039= i_window.window_13[02];
assign PB_039= i_window.window_17[07];
assign PA_040= i_window.window_13[12];
assign PB_040= i_window.window_18[13];
assign PA_041= i_window.window_24[09];
assign PB_041= i_window.window_06[11];
assign PA_042= i_window.window_27[23];
assign PB_042= i_window.window_22[25];
assign PA_043= i_window.window_24[15];
assign PB_043= i_window.window_18[16];
assign PA_044= i_window.window_10[22];
assign PB_044= i_window.window_05[26];
assign PA_045= i_window.window_09[02];
assign PB_045= i_window.window_15[04];
assign PA_046= i_window.window_22[25];
assign PB_046= i_window.window_16[27];
assign PA_047= i_window.window_12[09];
assign PB_047= i_window.window_27[09];
assign PA_048= i_window.window_06[25];
assign PB_048= i_window.window_11[27];
assign PA_049= i_window.window_23[02];
assign PB_049= i_window.window_03[07];
assign PA_050= i_window.window_15[02];
assign PB_050= i_window.window_11[07];
assign PA_051= i_window.window_18[18];
assign PB_051= i_window.window_23[22];
assign PA_052= i_window.window_22[20];
assign PB_052= i_window.window_08[25];
assign PA_053= i_window.window_22[14];
assign PB_053= i_window.window_03[16];
assign PA_054= i_window.window_05[18];
assign PB_054= i_window.window_21[20];
assign PA_055= i_window.window_11[17];
assign PB_055= i_window.window_05[18];
assign PA_056= i_window.window_15[02];
assign PB_056= i_window.window_20[02];
assign PA_057= i_window.window_08[02];
assign PB_057= i_window.window_27[03];
assign PA_058= i_window.window_18[02];
assign PB_058= i_window.window_23[04];
assign PA_059= i_window.window_27[08];
assign PB_059= i_window.window_22[11];
assign PA_060= i_window.window_05[21];
assign PB_060= i_window.window_23[27];
assign PA_061= i_window.window_14[06];
assign PB_061= i_window.window_09[08];
assign PA_062= i_window.window_10[13];
assign PB_062= i_window.window_27[15];
assign PA_063= i_window.window_20[03];
assign PB_063= i_window.window_20[08];
assign PA_064= i_window.window_05[18];
assign PB_064= i_window.window_02[23];
assign PA_065= i_window.window_08[08];
assign PB_065= i_window.window_20[11];
assign PA_066= i_window.window_13[12];
assign PB_066= i_window.window_08[14];
assign PA_067= i_window.window_24[17];
assign PB_067= i_window.window_04[20];
assign PA_068= i_window.window_02[04];
assign PB_068= i_window.window_02[10];
assign PA_069= i_window.window_21[14];
assign PB_069= i_window.window_14[15];
assign PA_070= i_window.window_12[20];
assign PB_070= i_window.window_17[20];
assign PA_071= i_window.window_02[11];
assign PB_071= i_window.window_27[11];
assign PA_072= i_window.window_09[06];
assign PB_072= i_window.window_21[06];
assign PA_073= i_window.window_05[03];
assign PB_073= i_window.window_11[07];
assign PA_074= i_window.window_17[25];
assign PB_074= i_window.window_12[27];
assign PA_075= i_window.window_27[22];
assign PB_075= i_window.window_27[27];
assign PA_076= i_window.window_02[08];
assign PB_076= i_window.window_20[09];
assign PA_077= i_window.window_24[11];
assign PB_077= i_window.window_19[12];
assign PA_078= i_window.window_14[22];
assign PB_078= i_window.window_17[27];
assign PA_079= i_window.window_21[08];
assign PB_079= i_window.window_16[10];
assign PA_080= i_window.window_26[02];
assign PB_080= i_window.window_20[03];
assign PA_081= i_window.window_22[12];
assign PB_081= i_window.window_09[13];
assign PA_082= i_window.window_07[22];
assign PB_082= i_window.window_08[27];
assign PA_083= i_window.window_08[02];
assign PB_083= i_window.window_03[04];
assign PA_084= i_window.window_12[16];
assign PB_084= i_window.window_27[27];
assign PA_085= i_window.window_09[17];
assign PB_085= i_window.window_15[18];
assign PA_086= i_window.window_18[11];
assign PB_086= i_window.window_02[13];
assign PA_087= i_window.window_02[14];
assign PB_087= i_window.window_24[16];
assign PA_088= i_window.window_16[22];
assign PB_088= i_window.window_09[23];
assign PA_089= i_window.window_14[16];
assign PB_089= i_window.window_27[18];
assign PA_090= i_window.window_16[24];
assign PB_090= i_window.window_21[27];
assign PA_091= i_window.window_06[14];
assign PB_091= i_window.window_18[14];
assign PA_092= i_window.window_02[02];
assign PB_092= i_window.window_20[05];
assign PA_093= i_window.window_22[22];
assign PB_093= i_window.window_27[25];
assign PA_094= i_window.window_10[27];
assign PB_094= i_window.window_24[27];
assign PA_095= i_window.window_18[21];
assign PB_095= i_window.window_26[22];
assign PA_096= i_window.window_02[20];
assign PB_096= i_window.window_25[21];
assign PA_097= i_window.window_03[17];
assign PB_097= i_window.window_18[17];
assign PA_098= i_window.window_23[18];
assign PB_098= i_window.window_09[19];
assign PA_099= i_window.window_21[17];
assign PB_099= i_window.window_02[27];
assign PA_100= i_window.window_03[24];
assign PB_100= i_window.window_18[25];
assign PA_101= i_window.window_19[07];
assign PB_101= i_window.window_24[08];
assign PA_102= i_window.window_27[04];
assign PB_102= i_window.window_09[11];
assign PA_103= i_window.window_27[16];
assign PB_103= i_window.window_07[17];
assign PA_104= i_window.window_06[21];
assign PB_104= i_window.window_11[22];
assign PA_105= i_window.window_18[17];
assign PB_105= i_window.window_13[18];
assign PA_106= i_window.window_18[21];
assign PB_106= i_window.window_15[26];
assign PA_107= i_window.window_12[18];
assign PB_107= i_window.window_07[23];
assign PA_108= i_window.window_23[22];
assign PB_108= i_window.window_18[24];
assign PA_109= i_window.window_10[04];
assign PB_109= i_window.window_11[09];
assign PA_110= i_window.window_26[05];
assign PB_110= i_window.window_25[10];
assign PA_111= i_window.window_07[10];
assign PB_111= i_window.window_27[12];
assign PA_112= i_window.window_20[05];
assign PB_112= i_window.window_15[06];
assign PA_113= i_window.window_14[23];
assign PB_113= i_window.window_09[27];
assign PA_114= i_window.window_09[19];
assign PB_114= i_window.window_04[21];
assign PA_115= i_window.window_27[05];
assign PB_115= i_window.window_22[07];
assign PA_116= i_window.window_13[19];
assign PB_116= i_window.window_22[21];
assign PA_117= i_window.window_15[13];
assign PB_117= i_window.window_27[13];
assign PA_118= i_window.window_07[10];
assign PB_118= i_window.window_17[10];
assign PA_119= i_window.window_09[22];
assign PB_119= i_window.window_27[25];
assign PA_120= i_window.window_02[06];
assign PB_120= i_window.window_07[07];
assign PA_121= i_window.window_02[10];
assign PB_121= i_window.window_13[10];
assign PA_122= i_window.window_07[23];
assign PB_122= i_window.window_02[24];
assign PA_123= i_window.window_04[06];
assign PB_123= i_window.window_15[06];
assign PA_124= i_window.window_07[16];
assign PB_124= i_window.window_13[16];
assign PA_125= i_window.window_11[22];
assign PB_125= i_window.window_16[24];
assign PA_126= i_window.window_16[13];
assign PB_126= i_window.window_11[14];
assign PA_127= i_window.window_09[26];
assign PB_127= i_window.window_04[27];
assign PA_128= i_window.window_06[03];
assign PB_128= i_window.window_19[09];
assign PA_129= i_window.window_22[18];
assign PB_129= i_window.window_27[22];
assign PA_130= i_window.window_20[20];
assign PB_130= i_window.window_23[25];
assign PA_131= i_window.window_11[15];
assign PB_131= i_window.window_23[17];
assign PA_132= i_window.window_27[06];
assign PB_132= i_window.window_02[10];
assign PA_133= i_window.window_22[15];
assign PB_133= i_window.window_27[17];
assign PA_134= i_window.window_17[14];
assign PB_134= i_window.window_22[16];
assign PA_135= i_window.window_26[20];
assign PB_135= i_window.window_06[22];
assign PA_136= i_window.window_20[18];
assign PB_136= i_window.window_07[21];
assign PA_137= i_window.window_11[02];
assign PB_137= i_window.window_24[07];
assign PA_138= i_window.window_24[10];
assign PB_138= i_window.window_12[12];
assign PA_139= i_window.window_08[11];
assign PB_139= i_window.window_03[12];
assign PA_140= i_window.window_20[21];
assign PB_140= i_window.window_15[23];
assign PA_141= i_window.window_21[08];
assign PB_141= i_window.window_27[09];
assign PA_142= i_window.window_21[02];
assign PB_142= i_window.window_13[10];
assign PA_143= i_window.window_05[16];
assign PB_143= i_window.window_25[18];
assign PA_144= i_window.window_16[19];
assign PB_144= i_window.window_11[23];
assign PA_145= i_window.window_13[13];
assign PB_145= i_window.window_02[17];
assign PA_146= i_window.window_03[17];
assign PB_146= i_window.window_27[27];
assign PA_147= i_window.window_02[13];
assign PB_147= i_window.window_09[15];
assign PA_148= i_window.window_16[19];
assign PB_148= i_window.window_18[24];
assign PA_149= i_window.window_05[09];
assign PB_149= i_window.window_10[12];
assign PA_150= i_window.window_02[12];
assign PB_150= i_window.window_16[14];
assign PA_151= i_window.window_20[22];
assign PB_151= i_window.window_04[27];
assign PA_152= i_window.window_13[19];
assign PB_152= i_window.window_08[20];
assign PA_153= i_window.window_24[02];
assign PB_153= i_window.window_10[06];
assign PA_154= i_window.window_16[22];
assign PB_154= i_window.window_21[23];
assign PA_155= i_window.window_07[22];
assign PB_155= i_window.window_21[22];
assign PA_156= i_window.window_11[08];
assign PB_156= i_window.window_16[08];
assign PA_157= i_window.window_26[07];
assign PB_157= i_window.window_07[08];
assign PA_158= i_window.window_21[02];
assign PB_158= i_window.window_07[03];
assign PA_159= i_window.window_19[17];
assign PB_159= i_window.window_24[18];
assign PA_160= i_window.window_10[25];
assign PB_160= i_window.window_18[27];
assign PA_161= i_window.window_10[09];
assign PB_161= i_window.window_22[09];
assign PA_162= i_window.window_12[23];
assign PB_162= i_window.window_07[24];
assign PA_163= i_window.window_03[17];
assign PB_163= i_window.window_23[17];
assign PA_164= i_window.window_13[04];
assign PB_164= i_window.window_18[05];
assign PA_165= i_window.window_02[03];
assign PB_165= i_window.window_06[08];
assign PA_166= i_window.window_15[04];
assign PB_166= i_window.window_10[05];
assign PA_167= i_window.window_12[20];
assign PB_167= i_window.window_23[26];
assign PA_168= i_window.window_02[13];
assign PB_168= i_window.window_27[14];
assign PA_169= i_window.window_07[14];
assign PB_169= i_window.window_24[15];
assign PA_170= i_window.window_04[02];
assign PB_170= i_window.window_10[03];
assign PA_171= i_window.window_13[05];
assign PB_171= i_window.window_26[05];
assign PA_172= i_window.window_24[12];
assign PB_172= i_window.window_02[13];
assign PA_173= i_window.window_12[17];
assign PB_173= i_window.window_17[18];
assign PA_174= i_window.window_02[06];
assign PB_174= i_window.window_15[11];
assign PA_175= i_window.window_21[11];
assign PB_175= i_window.window_05[12];
assign PA_176= i_window.window_27[11];
assign PB_176= i_window.window_08[13];
assign PA_177= i_window.window_04[09];
assign PB_177= i_window.window_24[11];
assign PA_178= i_window.window_12[21];
assign PB_178= i_window.window_26[21];
assign PA_179= i_window.window_26[02];
assign PB_179= i_window.window_20[10];
assign PA_180= i_window.window_26[26];
assign PB_180= i_window.window_21[27];
assign PA_181= i_window.window_10[22];
assign PB_181= i_window.window_13[27];
assign PA_182= i_window.window_27[14];
assign PB_182= i_window.window_22[15];
assign PA_183= i_window.window_07[11];
assign PB_183= i_window.window_13[12];
assign PA_184= i_window.window_16[08];
assign PB_184= i_window.window_22[09];
assign PA_185= i_window.window_03[02];
assign PB_185= i_window.window_02[07];
assign PA_186= i_window.window_13[08];
assign PB_186= i_window.window_07[09];
assign PA_187= i_window.window_20[07];
assign PB_187= i_window.window_06[09];
assign PA_188= i_window.window_14[10];
assign PB_188= i_window.window_20[11];
assign PA_189= i_window.window_22[02];
assign PB_189= i_window.window_25[07];
assign PA_190= i_window.window_20[16];
assign PB_190= i_window.window_02[20];
assign PA_191= i_window.window_15[16];
assign PB_191= i_window.window_02[25];
assign PA_192= i_window.window_27[24];
assign PB_192= i_window.window_14[25];
assign PA_193= i_window.window_07[20];
assign PB_193= i_window.window_06[25];
assign PA_194= i_window.window_26[14];
assign PB_194= i_window.window_02[16];
assign PA_195= i_window.window_12[06];
assign PB_195= i_window.window_17[09];
assign PA_196= i_window.window_05[14];
assign PB_196= i_window.window_27[16];
assign PA_197= i_window.window_16[02];
assign PB_197= i_window.window_05[07];
assign PA_198= i_window.window_04[23];
assign PB_198= i_window.window_09[25];
assign PA_199= i_window.window_02[17];
assign PB_199= i_window.window_09[18];
assign PA_200= i_window.window_02[22];
assign PB_200= i_window.window_06[27];
assign PA_201= i_window.window_05[05];
assign PB_201= i_window.window_08[10];
assign PA_202= i_window.window_07[05];
assign PB_202= i_window.window_02[07];
assign PA_203= i_window.window_09[19];
assign PB_203= i_window.window_20[23];
assign PA_204= i_window.window_27[18];
assign PB_204= i_window.window_02[23];
assign PA_205= i_window.window_17[11];
assign PB_205= i_window.window_12[12];
assign PA_206= i_window.window_02[20];
assign PB_206= i_window.window_03[25];
assign PA_207= i_window.window_02[19];
assign PB_207= i_window.window_14[20];
assign PA_208= i_window.window_24[06];
assign PB_208= i_window.window_18[11];
assign PA_209= i_window.window_18[15];
assign PB_209= i_window.window_06[18];
assign PA_210= i_window.window_16[03];
assign PB_210= i_window.window_16[09];
assign PA_211= i_window.window_17[18];
assign PB_211= i_window.window_07[19];
assign PA_212= i_window.window_05[05];
assign PB_212= i_window.window_24[05];
assign PA_213= i_window.window_02[23];
assign PB_213= i_window.window_27[27];
assign PA_214= i_window.window_03[07];
assign PB_214= i_window.window_10[09];
assign PA_215= i_window.window_17[17];
assign PB_215= i_window.window_22[18];
assign PA_216= i_window.window_21[25];
assign PB_216= i_window.window_07[26];
assign PA_217= i_window.window_23[21];
assign PB_217= i_window.window_03[23];
assign PA_218= i_window.window_25[08];
assign PB_218= i_window.window_20[09];
assign PA_219= i_window.window_06[12];
assign PB_219= i_window.window_24[12];
assign PA_220= i_window.window_02[14];
assign PB_220= i_window.window_20[14];
assign PA_221= i_window.window_08[12];
assign PB_221= i_window.window_19[12];
assign PA_222= i_window.window_13[07];
assign PB_222= i_window.window_18[07];
assign PA_223= i_window.window_17[19];
assign PB_223= i_window.window_27[27];
assign PA_224= i_window.window_10[17];
assign PB_224= i_window.window_26[18];
assign PA_225= i_window.window_06[21];
assign PB_225= i_window.window_02[26];
assign PA_226= i_window.window_14[18];
assign PB_226= i_window.window_27[22];
assign PA_227= i_window.window_14[26];
assign PB_227= i_window.window_19[27];
assign PA_228= i_window.window_15[12];
assign PB_228= i_window.window_21[12];
assign PA_229= i_window.window_04[19];
assign PB_229= i_window.window_27[19];
assign PA_230= i_window.window_11[17];
assign PB_230= i_window.window_16[17];
assign PA_231= i_window.window_09[05];
assign PB_231= i_window.window_16[07];
assign PA_232= i_window.window_22[02];
assign PB_232= i_window.window_16[04];
assign PA_233= i_window.window_27[02];
assign PB_233= i_window.window_02[04];
assign PA_234= i_window.window_15[21];
assign PB_234= i_window.window_02[26];
assign PA_235= i_window.window_14[15];
assign PB_235= i_window.window_19[16];
assign PA_236= i_window.window_18[02];
assign PB_236= i_window.window_13[06];
assign PA_237= i_window.window_23[06];
assign PB_237= i_window.window_12[09];
assign PA_238= i_window.window_09[02];
assign PB_238= i_window.window_13[07];
assign PA_239= i_window.window_06[20];
assign PB_239= i_window.window_25[23];
assign PA_240= i_window.window_22[17];
assign PB_240= i_window.window_06[18];
assign PA_241= i_window.window_09[14];
assign PB_241= i_window.window_14[14];
assign PA_242= i_window.window_20[24];
assign PB_242= i_window.window_13[26];
assign PA_243= i_window.window_12[26];
assign PB_243= i_window.window_07[27];
assign PA_244= i_window.window_15[18];
assign PB_244= i_window.window_20[18];
assign PA_245= i_window.window_19[14];
assign PB_245= i_window.window_25[15];
assign PA_246= i_window.window_09[18];
assign PB_246= i_window.window_20[19];
assign PA_247= i_window.window_15[02];
assign PB_247= i_window.window_20[05];
assign PA_248= i_window.window_23[20];
assign PB_248= i_window.window_26[27];
assign PA_249= i_window.window_24[23];
assign PB_249= i_window.window_09[24];
assign PA_250= i_window.window_11[22];
assign PB_250= i_window.window_03[23];
assign PA_251= i_window.window_19[05];
assign PB_251= i_window.window_24[05];
assign PA_252= i_window.window_18[22];
assign PB_252= i_window.window_19[27];
assign PA_253= i_window.window_08[24];
assign PB_253= i_window.window_13[25];
assign PA_254= i_window.window_15[22];
assign PB_254= i_window.window_13[27];
assign PA_255= i_window.window_09[14];
assign PB_255= i_window.window_04[15];


assign o_brief[000]=PA_000>PB_000 ? 1'b1 : 1'b0;
assign o_brief[001]=PA_001>PB_001 ? 1'b1 : 1'b0;
assign o_brief[002]=PA_002>PB_002 ? 1'b1 : 1'b0;
assign o_brief[003]=PA_003>PB_003 ? 1'b1 : 1'b0;
assign o_brief[004]=PA_004>PB_004 ? 1'b1 : 1'b0;
assign o_brief[005]=PA_005>PB_005 ? 1'b1 : 1'b0;
assign o_brief[006]=PA_006>PB_006 ? 1'b1 : 1'b0;
assign o_brief[007]=PA_007>PB_007 ? 1'b1 : 1'b0;
assign o_brief[008]=PA_008>PB_008 ? 1'b1 : 1'b0;
assign o_brief[009]=PA_009>PB_009 ? 1'b1 : 1'b0;
assign o_brief[010]=PA_010>PB_010 ? 1'b1 : 1'b0;
assign o_brief[011]=PA_011>PB_011 ? 1'b1 : 1'b0;
assign o_brief[012]=PA_012>PB_012 ? 1'b1 : 1'b0;
assign o_brief[013]=PA_013>PB_013 ? 1'b1 : 1'b0;
assign o_brief[014]=PA_014>PB_014 ? 1'b1 : 1'b0;
assign o_brief[015]=PA_015>PB_015 ? 1'b1 : 1'b0;
assign o_brief[016]=PA_016>PB_016 ? 1'b1 : 1'b0;
assign o_brief[017]=PA_017>PB_017 ? 1'b1 : 1'b0;
assign o_brief[018]=PA_018>PB_018 ? 1'b1 : 1'b0;
assign o_brief[019]=PA_019>PB_019 ? 1'b1 : 1'b0;
assign o_brief[020]=PA_020>PB_020 ? 1'b1 : 1'b0;
assign o_brief[021]=PA_021>PB_021 ? 1'b1 : 1'b0;
assign o_brief[022]=PA_022>PB_022 ? 1'b1 : 1'b0;
assign o_brief[023]=PA_023>PB_023 ? 1'b1 : 1'b0;
assign o_brief[024]=PA_024>PB_024 ? 1'b1 : 1'b0;
assign o_brief[025]=PA_025>PB_025 ? 1'b1 : 1'b0;
assign o_brief[026]=PA_026>PB_026 ? 1'b1 : 1'b0;
assign o_brief[027]=PA_027>PB_027 ? 1'b1 : 1'b0;
assign o_brief[028]=PA_028>PB_028 ? 1'b1 : 1'b0;
assign o_brief[029]=PA_029>PB_029 ? 1'b1 : 1'b0;
assign o_brief[030]=PA_030>PB_030 ? 1'b1 : 1'b0;
assign o_brief[031]=PA_031>PB_031 ? 1'b1 : 1'b0;
assign o_brief[032]=PA_032>PB_032 ? 1'b1 : 1'b0;
assign o_brief[033]=PA_033>PB_033 ? 1'b1 : 1'b0;
assign o_brief[034]=PA_034>PB_034 ? 1'b1 : 1'b0;
assign o_brief[035]=PA_035>PB_035 ? 1'b1 : 1'b0;
assign o_brief[036]=PA_036>PB_036 ? 1'b1 : 1'b0;
assign o_brief[037]=PA_037>PB_037 ? 1'b1 : 1'b0;
assign o_brief[038]=PA_038>PB_038 ? 1'b1 : 1'b0;
assign o_brief[039]=PA_039>PB_039 ? 1'b1 : 1'b0;
assign o_brief[040]=PA_040>PB_040 ? 1'b1 : 1'b0;
assign o_brief[041]=PA_041>PB_041 ? 1'b1 : 1'b0;
assign o_brief[042]=PA_042>PB_042 ? 1'b1 : 1'b0;
assign o_brief[043]=PA_043>PB_043 ? 1'b1 : 1'b0;
assign o_brief[044]=PA_044>PB_044 ? 1'b1 : 1'b0;
assign o_brief[045]=PA_045>PB_045 ? 1'b1 : 1'b0;
assign o_brief[046]=PA_046>PB_046 ? 1'b1 : 1'b0;
assign o_brief[047]=PA_047>PB_047 ? 1'b1 : 1'b0;
assign o_brief[048]=PA_048>PB_048 ? 1'b1 : 1'b0;
assign o_brief[049]=PA_049>PB_049 ? 1'b1 : 1'b0;
assign o_brief[050]=PA_050>PB_050 ? 1'b1 : 1'b0;
assign o_brief[051]=PA_051>PB_051 ? 1'b1 : 1'b0;
assign o_brief[052]=PA_052>PB_052 ? 1'b1 : 1'b0;
assign o_brief[053]=PA_053>PB_053 ? 1'b1 : 1'b0;
assign o_brief[054]=PA_054>PB_054 ? 1'b1 : 1'b0;
assign o_brief[055]=PA_055>PB_055 ? 1'b1 : 1'b0;
assign o_brief[056]=PA_056>PB_056 ? 1'b1 : 1'b0;
assign o_brief[057]=PA_057>PB_057 ? 1'b1 : 1'b0;
assign o_brief[058]=PA_058>PB_058 ? 1'b1 : 1'b0;
assign o_brief[059]=PA_059>PB_059 ? 1'b1 : 1'b0;
assign o_brief[060]=PA_060>PB_060 ? 1'b1 : 1'b0;
assign o_brief[061]=PA_061>PB_061 ? 1'b1 : 1'b0;
assign o_brief[062]=PA_062>PB_062 ? 1'b1 : 1'b0;
assign o_brief[063]=PA_063>PB_063 ? 1'b1 : 1'b0;
assign o_brief[064]=PA_064>PB_064 ? 1'b1 : 1'b0;
assign o_brief[065]=PA_065>PB_065 ? 1'b1 : 1'b0;
assign o_brief[066]=PA_066>PB_066 ? 1'b1 : 1'b0;
assign o_brief[067]=PA_067>PB_067 ? 1'b1 : 1'b0;
assign o_brief[068]=PA_068>PB_068 ? 1'b1 : 1'b0;
assign o_brief[069]=PA_069>PB_069 ? 1'b1 : 1'b0;
assign o_brief[070]=PA_070>PB_070 ? 1'b1 : 1'b0;
assign o_brief[071]=PA_071>PB_071 ? 1'b1 : 1'b0;
assign o_brief[072]=PA_072>PB_072 ? 1'b1 : 1'b0;
assign o_brief[073]=PA_073>PB_073 ? 1'b1 : 1'b0;
assign o_brief[074]=PA_074>PB_074 ? 1'b1 : 1'b0;
assign o_brief[075]=PA_075>PB_075 ? 1'b1 : 1'b0;
assign o_brief[076]=PA_076>PB_076 ? 1'b1 : 1'b0;
assign o_brief[077]=PA_077>PB_077 ? 1'b1 : 1'b0;
assign o_brief[078]=PA_078>PB_078 ? 1'b1 : 1'b0;
assign o_brief[079]=PA_079>PB_079 ? 1'b1 : 1'b0;
assign o_brief[080]=PA_080>PB_080 ? 1'b1 : 1'b0;
assign o_brief[081]=PA_081>PB_081 ? 1'b1 : 1'b0;
assign o_brief[082]=PA_082>PB_082 ? 1'b1 : 1'b0;
assign o_brief[083]=PA_083>PB_083 ? 1'b1 : 1'b0;
assign o_brief[084]=PA_084>PB_084 ? 1'b1 : 1'b0;
assign o_brief[085]=PA_085>PB_085 ? 1'b1 : 1'b0;
assign o_brief[086]=PA_086>PB_086 ? 1'b1 : 1'b0;
assign o_brief[087]=PA_087>PB_087 ? 1'b1 : 1'b0;
assign o_brief[088]=PA_088>PB_088 ? 1'b1 : 1'b0;
assign o_brief[089]=PA_089>PB_089 ? 1'b1 : 1'b0;
assign o_brief[090]=PA_090>PB_090 ? 1'b1 : 1'b0;
assign o_brief[091]=PA_091>PB_091 ? 1'b1 : 1'b0;
assign o_brief[092]=PA_092>PB_092 ? 1'b1 : 1'b0;
assign o_brief[093]=PA_093>PB_093 ? 1'b1 : 1'b0;
assign o_brief[094]=PA_094>PB_094 ? 1'b1 : 1'b0;
assign o_brief[095]=PA_095>PB_095 ? 1'b1 : 1'b0;
assign o_brief[096]=PA_096>PB_096 ? 1'b1 : 1'b0;
assign o_brief[097]=PA_097>PB_097 ? 1'b1 : 1'b0;
assign o_brief[098]=PA_098>PB_098 ? 1'b1 : 1'b0;
assign o_brief[099]=PA_099>PB_099 ? 1'b1 : 1'b0;
assign o_brief[100]=PA_100>PB_100 ? 1'b1 : 1'b0;
assign o_brief[101]=PA_101>PB_101 ? 1'b1 : 1'b0;
assign o_brief[102]=PA_102>PB_102 ? 1'b1 : 1'b0;
assign o_brief[103]=PA_103>PB_103 ? 1'b1 : 1'b0;
assign o_brief[104]=PA_104>PB_104 ? 1'b1 : 1'b0;
assign o_brief[105]=PA_105>PB_105 ? 1'b1 : 1'b0;
assign o_brief[106]=PA_106>PB_106 ? 1'b1 : 1'b0;
assign o_brief[107]=PA_107>PB_107 ? 1'b1 : 1'b0;
assign o_brief[108]=PA_108>PB_108 ? 1'b1 : 1'b0;
assign o_brief[109]=PA_109>PB_109 ? 1'b1 : 1'b0;
assign o_brief[110]=PA_110>PB_110 ? 1'b1 : 1'b0;
assign o_brief[111]=PA_111>PB_111 ? 1'b1 : 1'b0;
assign o_brief[112]=PA_112>PB_112 ? 1'b1 : 1'b0;
assign o_brief[113]=PA_113>PB_113 ? 1'b1 : 1'b0;
assign o_brief[114]=PA_114>PB_114 ? 1'b1 : 1'b0;
assign o_brief[115]=PA_115>PB_115 ? 1'b1 : 1'b0;
assign o_brief[116]=PA_116>PB_116 ? 1'b1 : 1'b0;
assign o_brief[117]=PA_117>PB_117 ? 1'b1 : 1'b0;
assign o_brief[118]=PA_118>PB_118 ? 1'b1 : 1'b0;
assign o_brief[119]=PA_119>PB_119 ? 1'b1 : 1'b0;
assign o_brief[120]=PA_120>PB_120 ? 1'b1 : 1'b0;
assign o_brief[121]=PA_121>PB_121 ? 1'b1 : 1'b0;
assign o_brief[122]=PA_122>PB_122 ? 1'b1 : 1'b0;
assign o_brief[123]=PA_123>PB_123 ? 1'b1 : 1'b0;
assign o_brief[124]=PA_124>PB_124 ? 1'b1 : 1'b0;
assign o_brief[125]=PA_125>PB_125 ? 1'b1 : 1'b0;
assign o_brief[126]=PA_126>PB_126 ? 1'b1 : 1'b0;
assign o_brief[127]=PA_127>PB_127 ? 1'b1 : 1'b0;
assign o_brief[128]=PA_128>PB_128 ? 1'b1 : 1'b0;
assign o_brief[129]=PA_129>PB_129 ? 1'b1 : 1'b0;
assign o_brief[130]=PA_130>PB_130 ? 1'b1 : 1'b0;
assign o_brief[131]=PA_131>PB_131 ? 1'b1 : 1'b0;
assign o_brief[132]=PA_132>PB_132 ? 1'b1 : 1'b0;
assign o_brief[133]=PA_133>PB_133 ? 1'b1 : 1'b0;
assign o_brief[134]=PA_134>PB_134 ? 1'b1 : 1'b0;
assign o_brief[135]=PA_135>PB_135 ? 1'b1 : 1'b0;
assign o_brief[136]=PA_136>PB_136 ? 1'b1 : 1'b0;
assign o_brief[137]=PA_137>PB_137 ? 1'b1 : 1'b0;
assign o_brief[138]=PA_138>PB_138 ? 1'b1 : 1'b0;
assign o_brief[139]=PA_139>PB_139 ? 1'b1 : 1'b0;
assign o_brief[140]=PA_140>PB_140 ? 1'b1 : 1'b0;
assign o_brief[141]=PA_141>PB_141 ? 1'b1 : 1'b0;
assign o_brief[142]=PA_142>PB_142 ? 1'b1 : 1'b0;
assign o_brief[143]=PA_143>PB_143 ? 1'b1 : 1'b0;
assign o_brief[144]=PA_144>PB_144 ? 1'b1 : 1'b0;
assign o_brief[145]=PA_145>PB_145 ? 1'b1 : 1'b0;
assign o_brief[146]=PA_146>PB_146 ? 1'b1 : 1'b0;
assign o_brief[147]=PA_147>PB_147 ? 1'b1 : 1'b0;
assign o_brief[148]=PA_148>PB_148 ? 1'b1 : 1'b0;
assign o_brief[149]=PA_149>PB_149 ? 1'b1 : 1'b0;
assign o_brief[150]=PA_150>PB_150 ? 1'b1 : 1'b0;
assign o_brief[151]=PA_151>PB_151 ? 1'b1 : 1'b0;
assign o_brief[152]=PA_152>PB_152 ? 1'b1 : 1'b0;
assign o_brief[153]=PA_153>PB_153 ? 1'b1 : 1'b0;
assign o_brief[154]=PA_154>PB_154 ? 1'b1 : 1'b0;
assign o_brief[155]=PA_155>PB_155 ? 1'b1 : 1'b0;
assign o_brief[156]=PA_156>PB_156 ? 1'b1 : 1'b0;
assign o_brief[157]=PA_157>PB_157 ? 1'b1 : 1'b0;
assign o_brief[158]=PA_158>PB_158 ? 1'b1 : 1'b0;
assign o_brief[159]=PA_159>PB_159 ? 1'b1 : 1'b0;
assign o_brief[160]=PA_160>PB_160 ? 1'b1 : 1'b0;
assign o_brief[161]=PA_161>PB_161 ? 1'b1 : 1'b0;
assign o_brief[162]=PA_162>PB_162 ? 1'b1 : 1'b0;
assign o_brief[163]=PA_163>PB_163 ? 1'b1 : 1'b0;
assign o_brief[164]=PA_164>PB_164 ? 1'b1 : 1'b0;
assign o_brief[165]=PA_165>PB_165 ? 1'b1 : 1'b0;
assign o_brief[166]=PA_166>PB_166 ? 1'b1 : 1'b0;
assign o_brief[167]=PA_167>PB_167 ? 1'b1 : 1'b0;
assign o_brief[168]=PA_168>PB_168 ? 1'b1 : 1'b0;
assign o_brief[169]=PA_169>PB_169 ? 1'b1 : 1'b0;
assign o_brief[170]=PA_170>PB_170 ? 1'b1 : 1'b0;
assign o_brief[171]=PA_171>PB_171 ? 1'b1 : 1'b0;
assign o_brief[172]=PA_172>PB_172 ? 1'b1 : 1'b0;
assign o_brief[173]=PA_173>PB_173 ? 1'b1 : 1'b0;
assign o_brief[174]=PA_174>PB_174 ? 1'b1 : 1'b0;
assign o_brief[175]=PA_175>PB_175 ? 1'b1 : 1'b0;
assign o_brief[176]=PA_176>PB_176 ? 1'b1 : 1'b0;
assign o_brief[177]=PA_177>PB_177 ? 1'b1 : 1'b0;
assign o_brief[178]=PA_178>PB_178 ? 1'b1 : 1'b0;
assign o_brief[179]=PA_179>PB_179 ? 1'b1 : 1'b0;
assign o_brief[180]=PA_180>PB_180 ? 1'b1 : 1'b0;
assign o_brief[181]=PA_181>PB_181 ? 1'b1 : 1'b0;
assign o_brief[182]=PA_182>PB_182 ? 1'b1 : 1'b0;
assign o_brief[183]=PA_183>PB_183 ? 1'b1 : 1'b0;
assign o_brief[184]=PA_184>PB_184 ? 1'b1 : 1'b0;
assign o_brief[185]=PA_185>PB_185 ? 1'b1 : 1'b0;
assign o_brief[186]=PA_186>PB_186 ? 1'b1 : 1'b0;
assign o_brief[187]=PA_187>PB_187 ? 1'b1 : 1'b0;
assign o_brief[188]=PA_188>PB_188 ? 1'b1 : 1'b0;
assign o_brief[189]=PA_189>PB_189 ? 1'b1 : 1'b0;
assign o_brief[190]=PA_190>PB_190 ? 1'b1 : 1'b0;
assign o_brief[191]=PA_191>PB_191 ? 1'b1 : 1'b0;
assign o_brief[192]=PA_192>PB_192 ? 1'b1 : 1'b0;
assign o_brief[193]=PA_193>PB_193 ? 1'b1 : 1'b0;
assign o_brief[194]=PA_194>PB_194 ? 1'b1 : 1'b0;
assign o_brief[195]=PA_195>PB_195 ? 1'b1 : 1'b0;
assign o_brief[196]=PA_196>PB_196 ? 1'b1 : 1'b0;
assign o_brief[197]=PA_197>PB_197 ? 1'b1 : 1'b0;
assign o_brief[198]=PA_198>PB_198 ? 1'b1 : 1'b0;
assign o_brief[199]=PA_199>PB_199 ? 1'b1 : 1'b0;
assign o_brief[200]=PA_200>PB_200 ? 1'b1 : 1'b0;
assign o_brief[201]=PA_201>PB_201 ? 1'b1 : 1'b0;
assign o_brief[202]=PA_202>PB_202 ? 1'b1 : 1'b0;
assign o_brief[203]=PA_203>PB_203 ? 1'b1 : 1'b0;
assign o_brief[204]=PA_204>PB_204 ? 1'b1 : 1'b0;
assign o_brief[205]=PA_205>PB_205 ? 1'b1 : 1'b0;
assign o_brief[206]=PA_206>PB_206 ? 1'b1 : 1'b0;
assign o_brief[207]=PA_207>PB_207 ? 1'b1 : 1'b0;
assign o_brief[208]=PA_208>PB_208 ? 1'b1 : 1'b0;
assign o_brief[209]=PA_209>PB_209 ? 1'b1 : 1'b0;
assign o_brief[210]=PA_210>PB_210 ? 1'b1 : 1'b0;
assign o_brief[211]=PA_211>PB_211 ? 1'b1 : 1'b0;
assign o_brief[212]=PA_212>PB_212 ? 1'b1 : 1'b0;
assign o_brief[213]=PA_213>PB_213 ? 1'b1 : 1'b0;
assign o_brief[214]=PA_214>PB_214 ? 1'b1 : 1'b0;
assign o_brief[215]=PA_215>PB_215 ? 1'b1 : 1'b0;
assign o_brief[216]=PA_216>PB_216 ? 1'b1 : 1'b0;
assign o_brief[217]=PA_217>PB_217 ? 1'b1 : 1'b0;
assign o_brief[218]=PA_218>PB_218 ? 1'b1 : 1'b0;
assign o_brief[219]=PA_219>PB_219 ? 1'b1 : 1'b0;
assign o_brief[220]=PA_220>PB_220 ? 1'b1 : 1'b0;
assign o_brief[221]=PA_221>PB_221 ? 1'b1 : 1'b0;
assign o_brief[222]=PA_222>PB_222 ? 1'b1 : 1'b0;
assign o_brief[223]=PA_223>PB_223 ? 1'b1 : 1'b0;
assign o_brief[224]=PA_224>PB_224 ? 1'b1 : 1'b0;
assign o_brief[225]=PA_225>PB_225 ? 1'b1 : 1'b0;
assign o_brief[226]=PA_226>PB_226 ? 1'b1 : 1'b0;
assign o_brief[227]=PA_227>PB_227 ? 1'b1 : 1'b0;
assign o_brief[228]=PA_228>PB_228 ? 1'b1 : 1'b0;
assign o_brief[229]=PA_229>PB_229 ? 1'b1 : 1'b0;
assign o_brief[230]=PA_230>PB_230 ? 1'b1 : 1'b0;
assign o_brief[231]=PA_231>PB_231 ? 1'b1 : 1'b0;
assign o_brief[232]=PA_232>PB_232 ? 1'b1 : 1'b0;
assign o_brief[233]=PA_233>PB_233 ? 1'b1 : 1'b0;
assign o_brief[234]=PA_234>PB_234 ? 1'b1 : 1'b0;
assign o_brief[235]=PA_235>PB_235 ? 1'b1 : 1'b0;
assign o_brief[236]=PA_236>PB_236 ? 1'b1 : 1'b0;
assign o_brief[237]=PA_237>PB_237 ? 1'b1 : 1'b0;
assign o_brief[238]=PA_238>PB_238 ? 1'b1 : 1'b0;
assign o_brief[239]=PA_239>PB_239 ? 1'b1 : 1'b0;
assign o_brief[240]=PA_240>PB_240 ? 1'b1 : 1'b0;
assign o_brief[241]=PA_241>PB_241 ? 1'b1 : 1'b0;
assign o_brief[242]=PA_242>PB_242 ? 1'b1 : 1'b0;
assign o_brief[243]=PA_243>PB_243 ? 1'b1 : 1'b0;
assign o_brief[244]=PA_244>PB_244 ? 1'b1 : 1'b0;
assign o_brief[245]=PA_245>PB_245 ? 1'b1 : 1'b0;
assign o_brief[246]=PA_246>PB_246 ? 1'b1 : 1'b0;
assign o_brief[247]=PA_247>PB_247 ? 1'b1 : 1'b0;
assign o_brief[248]=PA_248>PB_248 ? 1'b1 : 1'b0;
assign o_brief[249]=PA_249>PB_249 ? 1'b1 : 1'b0;
assign o_brief[250]=PA_250>PB_250 ? 1'b1 : 1'b0;
assign o_brief[251]=PA_251>PB_251 ? 1'b1 : 1'b0;
assign o_brief[252]=PA_252>PB_252 ? 1'b1 : 1'b0;
assign o_brief[253]=PA_253>PB_253 ? 1'b1 : 1'b0;
assign o_brief[254]=PA_254>PB_254 ? 1'b1 : 1'b0;
assign o_brief[255]=PA_255>PB_255 ? 1'b1 : 1'b0;


endmodule