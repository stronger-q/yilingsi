`define IP_UUID _loopback_test                              
`define IP_NAME_CONCAT(a,b) a``b                            
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID) 
//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2023 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = efx_csi2_tx
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Tue May 30 16:05:37 2023
// ***************************************************************************************

`timescale 1 ns / 1 ps
module efx_csi2_tx_modelsim #(
    parameter tLPX_NS = 50,
    parameter tINIT_NS = 100000,
    parameter tINIT_SKEWCAL_NS = 100000,
    parameter tLP_EXIT_NS = 100,
    parameter tCLK_ZERO_NS = 262,
    parameter tCLK_TRAIL_NS = 60,
    parameter tCLK_POST_NS = 60,
    parameter tCLK_PRE_NS = 10,
    parameter tCLK_PREPARE_NS = 38,
    parameter tHS_PREPARE_NS = 40,
    parameter tWAKEUP_NS = 1000,
    parameter tHS_EXIT_NS = 100,
    parameter tHS_ZERO_NS = 105,
    parameter tHS_TRAIL_NS = 60,
    parameter NUM_DATA_LANE = 4,
    parameter HS_BYTECLK_MHZ = 100,
    parameter CLOCK_FREQ_MHZ = 100,
    parameter DPHY_CLOCK_MODE = "Continuous", 
    parameter PACK_TYPE = 4'b1111,
    parameter PIXEL_FIFO_DEPTH = 2048,  
    parameter ENABLE_VCX = 0,
    parameter FRAME_MODE = "GENERIC",    
    parameter ASYNC_STAGE = 2
)(
    input logic           reset_n,
    input logic           clk,				
    input logic           reset_byte_HS_n,
    input logic           clk_byte_HS,
    input logic           reset_pixel_n,
    input logic           clk_pixel,
	output logic          Tx_LP_CLK_P,
	output logic          Tx_LP_CLK_P_OE,
	output logic          Tx_LP_CLK_N,
	output logic          Tx_LP_CLK_N_OE,
	output logic [7:0]    Tx_HS_C,
	output logic          Tx_HS_enable_C,
    output logic [NUM_DATA_LANE-1:0]         Tx_LP_D_P,
    output logic [NUM_DATA_LANE-1:0]         Tx_LP_D_P_OE,
	output logic [NUM_DATA_LANE-1:0]         Tx_LP_D_N,
    output logic [NUM_DATA_LANE-1:0]         Tx_LP_D_N_OE,
	output logic [7:0]                       Tx_HS_D_0,
	output logic [7:0]                       Tx_HS_D_1,
	output logic [7:0]                       Tx_HS_D_2,
	output logic [7:0]                       Tx_HS_D_3,
	output logic [7:0]                       Tx_HS_D_4,
	output logic [7:0]                       Tx_HS_D_5,
	output logic [7:0]                       Tx_HS_D_6,
	output logic [7:0]                       Tx_HS_D_7,
	output logic [NUM_DATA_LANE-1:0]         Tx_HS_enable_D,
    input  logic          axi_clk,
    input  logic          axi_reset_n,
    input  logic   [5:0]  axi_awaddr,
    input  logic          axi_awvalid,
    output logic          axi_awready,
    input  logic   [31:0] axi_wdata,
    input  logic          axi_wvalid,
    output logic          axi_wready,
    output logic          axi_bvalid,
    input  logic          axi_bready,
    input  logic   [5:0]  axi_araddr,
    input  logic          axi_arvalid,
    output logic          axi_arready,
    output logic   [31:0] axi_rdata,
    output logic          axi_rvalid,
    input                 axi_rready,
    input logic           hsync_vc0,
    input logic           hsync_vc1,
    input logic           hsync_vc2,
    input logic           hsync_vc3,
    input logic           vsync_vc0,
    input logic           vsync_vc1,
    input logic           vsync_vc2,
    input logic           vsync_vc3,
    input logic           hsync_vc4,
    input logic           hsync_vc5,
    input logic           hsync_vc6,
    input logic           hsync_vc7,
    input logic           hsync_vc8,
    input logic           hsync_vc9,
    input logic           hsync_vc10,
    input logic           hsync_vc11,
    input logic           hsync_vc12,
    input logic           hsync_vc13,
    input logic           hsync_vc14,
    input logic           hsync_vc15,
    input logic           vsync_vc4,
    input logic           vsync_vc5,
    input logic           vsync_vc6,
    input logic           vsync_vc7,
    input logic           vsync_vc8,
    input logic           vsync_vc9,
    input logic           vsync_vc10,
    input logic           vsync_vc11,
    input logic           vsync_vc12,
    input logic           vsync_vc13,
    input logic           vsync_vc14,
    input logic           vsync_vc15,
    input logic [5:0]     datatype,   
    input logic [63:0]    pixel_data,
    input logic           pixel_data_valid,
    input logic [15:0]    haddr,   
    input logic [15:0]    line_num,
    input logic [15:0]    frame_num,
    output logic          irq
);
//pragma protect
//pragma protect begin
`protected

    MTI!#lU+ZJU}{Kos2B7mY#'sYx^_3=CO>W=,j"7Z[#=moCXG1$A$zsE\{pmsR$\KU2*oQE@E"k{w
    E5JvZw|'I!Tr!}O?l7GBG<v\e**ARYs}KuoRl3OK5le%L$}u1G^\=J-e^e*{V_><-RA<[X7BeQRk
    A'bJ[QUvCJp*[*=mBk~TEW]=X{R[DAYRN1#'K}ZGK|XUvO<[@T<+R]Q3JUZjvH@xXYo_3VEIj!z)
    \>3A2jBH]XnV7zi@<Ol$=R}I8E3*jJr3*Qw;=Y*G#-^EJQlmk@p@'w1Ejm^i,\7Z]TnV7WwwQks~
    ^.w^=o]R!el~!$HxD,@X3r_oU;^kW,XDe}hjIv1?1l}o1n?*C]im<D#-UKr#{-}+<VHo'>s1+B>w
    [[sB;&zOE>eW7OUa,e@s]u*zKXlsVR$]QET<RzRaxAc>>$v!XB2VkTYo@z2W1,55]u{H7{3la}$*
    U-<-T-Ip=BnExkuK7_E%}Ru,,3p;uSj}-<3v;QOKC#,Vu$Wzv<ct#DJDiX<n$SIv?C7Eor^2Z'T'
    Ars<5;D<>eFg'tcCZseR><#o7GGbS*{VsdC2T3GXaK]arTq?p5p!aKUw'=R=DWE1Sm+-+>$aB2Re
    u?U5-*8uAvY;H-ogixkDgxDZ71mVY9QUZ'v17Ag^Ozo^;GTE|\$G^S+ov#5-1{~AW[~{n-*{}"ju
    BIDIG>UCQQH_URjj+K,3>Ev5V_xk-_d]QBQ[#->}\'QRJYv_j^VDIZ-,Goul_'APZo3Y~<<XuYq\
    +{37?Gk[DnVfHn'!h:Aa]U-XaHlXjnOzYT,%+5#la^Du35,r5mza3Q?rI2oz(H[-VLD<T].FDs'a
    =eo}nU^-F'H$+\nTp-*!R>r?-YEl>R*1Ef,GXOZ5-VWjk[U{l~arll;Cmm3<z#IC5O$s'K^_I]~s
    ,A}3x2ljVK,;mBuD=vdCrKW2r1aBQQsX<YGsI+THX<<=e{mB*B'~rX~dQ]$*[-,{2Vk7r2G<+]pT
    <OZG6p"doK3?!e<]]C_ZI@z_^2T*Cl+3{=1]]~RZ7^>jRFIA{}le;;tq?[1EuBu;/>nA!?7oe)*!
    DwWCyQBDA6i7Ba^k'RxE1ZFHR#Cp7C3'rev_znUQ{5CU=[AYp;r]-e*RO-?w}kT#j?KGKVoSxmXI
    RG+apeln1GG2v\*^/@DKBoH_7]=x+'3Q>^0yA,,v*pD'=zI+r\YoYs>^m,Q-7}3*q*CwAAURikav
    \D{T<<5Ov^Zm1zW\z{$oGrZ@mQ#]vB5D-TQI*lHJ3H}G<#^$=N?<Q,p\]w_ilo)_KGw?VpHQ1{>Q
    [vmI[x5p#wO#EoDuajV~>AEk1nj:,}pBCs+wo,#2kIE$z'@-yIE]w{$x<j$DU)IBX~YmT{ei]xio
    jHTr@VG4#OU3{YTTm}Y?KTTC#<-3vD[?3{o#Ur!UA[1UvB#,R5x\as[k?UAKxvE7M_oXCQI#$w5B
    >=^V1p#K^}pGYRID^I3J=soe'3{VIRe>*=s>~GWUOa+R_xZeA{^}]D1wJI8'x{w!j+Tu=}Y1={7p
    ]+{{=\GKeUkK+o2QD2Q)f]D7sX=*mbe7QBuO,Kz~*<LPBK=Q,J<jYxBU9?GIG!VBrrAHjo>x{27C
    r2s;nR'u;8,A=j3^\C)EEY_eHsjIVkuCXn-<UDk%}+ZQ)~\[x=_lj<s<#jx-?+xGm/a*e[_UAo@I
    [x=oeD\+QZe'WVjI#v1!2!a\E!*B<?-]@YLi{BX[1iUR3YzoZGH.C=?of}ZQw-1+HRR_\KYVK$A$
    s;}]**Dv}iTujsZ!GThoam*?Esk{R5uXEUrl\DsnOpD|6E$inwU{z,$<,]_12\oZIOH;+xJ+s~<e
    CZNmV#^5knr~_XGvuHAIVY#JYR71Bn7-<R*\YY5oV'+>pYT['}U)p#wsR0sCnv$sO2z}J2dn=\*{
    I<3F-.XE-QnY2@BlUp\\1Y2'o7>{u2wA2pQssXEv3{UoAonHu{,p!sQU>peaW1Q,xeQYzk\#plHU
    ![u=keHIiU5!E1{Vm5C_p=1n<xIQlA;r3-Y?@!rv'${{Y;$z'1/E;+Cv5~u9pVVpKXHY0[#rY}we
    jBQ~Rx,YK\G;*R^,{almBl<p*6a,k\Dae+2Du'ioT3K>7GpzK>lu_v-x[QO}rkq#[_{K<T$?D^Wm
    sDAW,ax*TH~_s[Tis$Y\DTJ)PKov3ua$*Gu-2BIll}V<P8Yx{~1{XC,{pvW1u7ImI@vv-rl5}?XC
    #V'rv?Gx5m0gB\G~>z-}pX_]PRAWEbQYYV@pHw-p{@oTe]@TurYC_H9ruA!;BeEo^o~o-~Y112,2
    'A{;>j}x_jeEz5ux_1H;<U_Ope5bz_2^6@TeQAayD#>l=5VaOO1jP|_1WWY*>{1>J,_1BGsrw_1G
    ,{qsozIaG~'aR!IRm@<G7x2h_}w~5C>k:{&\D]\p'{]{'DR#<[X{T33'\7[%x^*~[3sEHo7]!oXx
    $lE#va;<f#Hrpd\B:I5VA^Ym5yn{ErvCspqW=wj5n}5\HVD[pDEE~ozY^oYssIRmEwrb1la_G}1@
    2\##~C5un-UWstBEvj2+ws7~Uk%GQxXa<O=^]7*gZQuOpzx~-GiJkUx>~Q]ew>>eBjvK-1'\0VB,
    3nz5!G-Aj}xppMT^_{^El=aIKRrR7zdOmRGr6nI5mk>^K_j]Jk,Ii#Vm1'!8a1I~=5lrk,r2$wla
    {'\AiXU_}Gu^>XaCB@!pvIkoxI@K=T>vh:QBI@Ik5JnDQZeXp[IY1?.1!R><rz7JrkJ;_TeY+w#T
    ]TAV}jJ/xJ5enzW}35lZjoTOWn$^K<}=^{I@TUDjABoIi=^G{TTv\VwB5eA;#+\VEE0P;>WwiDRl
    Wlsl5O;A~ll_^nEso|pHmU8251#D5aX}3jYUCH_9QZ^1zB^@pkCJyKo_'$T=l!U$@X>-CXU[xi'o
    @Y?O*OG2Ru{1e?oWapQYuZRv]G]{Yupe]~\Zm,GT!,7*23-,Te;['[kpJFzVe+Jw><R?_!XH3Q~X
    p5naZl^\H^=)r_*H*i!{x]-[*HG!67"17o,b/~XI]QCO]^CK+#5wT^K+o$,H[~Viz=dmx+{Ro>O!
    v7A}}k[in'n_an7
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#}a*prpDKvB*!RwvHaOa;x}W@WIoUURYW}Z-Wm&^i7@t~U=?^oWw[X^\0}0LwHACt}B{eU]i
    G-'@#[mlz77?@}aJ35/o_n=['CW!Ul$HUl=U7BvVO#oskU2*3vH!'#Z-C_Gs_KH9,@Ce|)v++ot1
    xl@r?jHNj;Xo]g}ZJQVK!?N5CD-^sz50)^Rm*^a,mx*R^uoB?\='E-DGK>&ov3^Z',?nl@av^l}Z
    DYm]{-X\!EHvA'^97$+n}m^A%}Vu[Y+RY!|KA^XQmRH$D-+<,G@fpz\$mo?pKYjr'zTuQ$i]Vmz@
    Di]\W&nj5!1x1CosorzxGDQzVs['[RzkTr.%i]V<uTK1-CYrS]'U#Ollre=2QBHmX$Kpuz[,H_$o
    AI7k@r^}k[~[no_o$W$oeRv!2lr<,NQuaQt?<p72EC{nO?CGWzlVW~e$+}UG;u<U-]Z]xk*q5zBU
    ujCzu_xZC[?;7#=YN+OW+[5?+o$m}_e]='1?5*kY'[O!pOT]u{w1Ai$W;;{-Z*\r~lQOpIapvYan
    [e\Xu37DWw<AZ5#+#$nMVQ{ZxZpWmY3*H-{IFVJ@o7*rVLij3j\_kwBV@a7+UlIO2WYnmQvX_~&A
    \W^@Xj<'pV3:J7l}B]i2o2Y~,ez^[Iwm(1,zi\7v\/Yg,BiC,roaNo}O,ACV$R$xE5Uw[L7^X\_@
    s^}jJaD;-u3a{7VZV![JO+BekGz*Cu4'DQ[$?jvOI7sjln-GKV,lGxu?Dl!;C-m$&={{E]!Q$JnE
    {QOgm]7Zf#^xoB]#m\eGs'^BaGZ'?IDM_VQHpquTX\ri\,#,e#%LQaneWz1^E5K^jUTow5Yk5s{I
    7#Jxw]]?=*+EAqKBr<pxaunjkX_nOD0*jkaDd\WVOIE$nYr5~]o7@ou=Z1zYnRVQ}l!),UCDT5<\
    |L8\[$J>EERK'!IIlC3l{@QN,3X!^~n_]l\ex]n]7WC[qixRij]>ATEp>?Ow#@T[Y>Uax,pE*BU]
    o!}ippx;!IZnV]aBx_,X<DW\e<^uJBTY@KzI3Hw>sv@HWZ1p}}p?@=elH=xnR><<J7+ppe2O{73*
    z@Dov@zReY+\!n>YIGz+w+[Tsu-@~qyajmesY2CRI*o,'#5TD#2?[g+-@eClKU'3aoqtx1{?R<+A
    [a]ef1U3;\<'}G><1^'''YX7*=IxzXxKzk_3*xuT^7?}]^-5rR5=pr3'VI1wXs?mVa1-;@X!562p
    QvMw\~<B>2T}x~Bq7Z<v}HYu1O_D~GQ3.c1T;~XX1~><Di^],]YxR3*5emOjUjO)~DooNJ{;<-l~
    ]Cm21?A>+HH{UC2aOs@z-iHIZ,{<Wz*A3VOORv^o,:lupi-Gl'k]R}iRi7SoCY!'m!1,Y[lB]EBB
    +5!:UX1@BA$YrG]@EB}3Ve*3r_X>T5lzUXI{Dk_17k_GI;slW{=Y@\C253OW#Te7CII2pIu[mRBk
    -5opazZpAv~usVnrs*Q7\n~H<l$]v~VK2jG7O,u!eH-H'uV^Y3+r3o3'ck\>R*us$lr_zaQ1u'+;
    p5<]T2>E^i=Q#I25<Q^GaljzRIm$rEE,Qi1-1e^DAvom5Zz+}[zIJo;_VTO\3,wKE]?QWIpwxLKD
    D_<'J#'[?w=+rotY>XZ[Zo,oDzn=D+^Ux3G=,]$o_Y_WDsDcr7p~sB<Zz<X7fT<m!}2,TkR~\j1O
    AEStl^[3Y=TKV5<3p>KEC#[zQv~Eo![^C@WY7[R+T{I>y;EaY2lEKiYZ@#eI{xE='CJ1@G5]pxK]
    #uz=HAxI;zBe#11$?avE5ix[z}vHx+=U'GvZo,35v[z'uX{mzaIIx\7R$QkAH=jV^vKIH)\DEkA[
    ?*Gl=XK+nou{5#m,l9rDXVrYKxEw+Hizz3~oz1f*uD!s!p'c;Bp}9:}[w1-=Irx7w22HQ5VI^V'B
    #owoC*$Hnu>'CzOnH1*iaYJ}IQEV;2VH5zsuYQIz{=B7QoX$2EsVm'5?TKr;[j13Ho^n$_aO7eVB
    'IA[,E+C7Yhz+QaC1D+Br@OWDE<V<5ZRT^?7J\<?YEkKn-TzCxTqb\{{\#T2>[)-}JrJw{aQxXBv
    Z}>ur;#]IY,?on[OumV@Cv<1[
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#j]vVuQ2;Ax1Xj1!Z|#w*Q'[il~Ya]lwb|%#&"[l}k>oUY!v3T<+Fv%2BmZIAW?jJRu7IaR-
    {AC@X=pgaap<+1$'Q,AmOoXA31,['>Kj^iY\|_j-RJ+z[v5Xe;TGR_$Cpek][omYK$@=ekU~p<*n
    '[+Ar;'$UreU,g=!x7aYQ*,O{I)eYH}eWx,=]1sZwjDzj#]K_jTkBrDI+<s>5*3rk-jpp\e5X<}{
    $#2[}'oJz'*$Qjr}'><Om,;i5oV'_?pupETO-Ojo'=x!,\*GlWssCD>Ba2zlsk?r*_i2XTk_'i1#
    sD*DH=Ook3_]#vC^2$$}_jiOiu>!+*luC~<I?XCCmmX<O-1Os2x_J~BQm{B}{ua*5kTz^}7#,1Uq
    [l\OIA[nzW'kzsVWTa@5p\HWC=\5S!sB,{YEm~$A2Je@$h=m'^arpkI'5@Rn->V>7-p'i59[?CBN
    1iKw1u{Kx>=j?]I3m7?l_*upgiwVDP{Y;!]e'Xg<<;BKaaKo<2}Nve$$2-$\'[$\!YRu!H,lV1ET
    1<BB|1;Ol=5e_7k]D'!pGHr~^^jaIYYioY5!uq?1?_?C*ITQBV_[rUUEYu*#eX}4Q=V{yuns@VR;
    a7uB?C7e5Le<
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#J[Z!>ez>1wnG-V<52vH,\Too{o'OH{>s}~{{p]#!Rr!]{7W*]'XDiHeI1'kr?5<$1-aEcY,
    Ham{_3N}mBz77?@}aJ35/o_n=['CW!Ul$HUl=U7BvVO#oskUm*3vH!'#Z-C_Gs_!H9,~CA|Q2pj]
    pQEVuX7;Hpij;Xo]g}ZJQVK!?N5CD-^sz5;QR=RWXG[vzRmsx'D@XeCW[!R1eGYmjm,jJC8Y#<T=
    Hji}ioWP>A_~}J'U*n~OHjUTi>K+gNi_pYz_{-*@B]JsvU5u<;5#2UGIwk7[3um}zm>1?sBmX;Z]
    3U;{rYeH0K{HH'g|=BBr*VrEi7X[x}kjwwvo>R2xBWrzva+OGr=$GQ;W_o7VcVzQDEa{rf\RUCa=
    K?pa\~x~\_Dj<A*w3a]--_]zp]/!=R7'[Je*-wXD_u=oYYGz4D!e_y9:K\sAmB!C/2(0Qc2Eu5&J
    GHlEYl^L~}wBv9oumjC7~]=!-7J=;+5H<sjzI297^$zHl=lUv?mGM[7,Wp3\{sDv==n[}]2[,=Zo
    kpk<a'RpaOjQRB>oIXoKuR#p~C$\m(w7W3,K~wDs#7iDu<6*}X{2ji<PB=D7UTQ<}lZYeo~]_oJ<
    ~,_oW$<>G@TQ<_r#z7_Rje!u+]r=2Q?^i8I[1B'~Eps2v>e,~Gc\/~]k~BzpX?p?G-su_Y\-+u}[
    VQ'w<<UI~5wVIQk!wQ[=eC^1uWw\osu^'DkpC{n}Q~aez:O-eW'lVn0uR^~7O~@<A$ZwUJmYY{~n
    +.IU{vtUI5w_THWuQk$EajK<>T^EW>KI,Z*k={IjzW+OkR_UDI*6[i_QC=eH?s@\13Q{KTx5Xe25
    }#K#vaDi3[Z*~eZRJA1WOeeH#n*~2-*?zOK=zuBs1KpZe~{*a,\xI;D_aUv+kT$^}"$C#>d>]Upm
    |v\}j$3DJu7W^xEU@K1[vmY@ZpAZjuE^[BVj\TwOO[k\>C~ZTri5@CbhJ5TY}i}@GOYa733BQoG{
    L#7m[TIi~-zW}eZO$$svYE<nKuw]Y#XO^xW-r)$<*-:+'rUinfm>@IF>o=l1I-kHe\@l_R>{]D<=
    RxlNlipvV1k@uB>X8Eo^Qjk}]pW~aE3T=1kB#Y_n+HRjYI?DC2BZ#sp,rC[;}hE~l$G_?Btsp][A
    5-7_zQ-T7J}$yVKC,Law11]5-5kGi7Ck!5Vj#Jmzra2zp>iaJ<i}kzzOYwe!2**Mlks5kpA!\#m$
    5J'lT<<n,<X74;E-'TQO"vx;r5~1-$!_1AR@ZjlZzGx<*1nD_Y'5mwj'7"p+J^B~O?@>;;,R>C%l
    XT3TUaui-Rw2-\@dI[<GfCCR*Kv;aH1-ah=iWl=T1I<lJREo?a&,E1otkOJK$Y3uRo[1UTo=W<J&
    Us+~j;]Wl@H3=OnJvz;I@D$s!n7udMx2VZkDD;rYnujZj>^[QZ2=v?dr3QI]GAr'5116?]XwI1@\
    DM*]7lz>3J(rv_,A{e!e{J>UaeIj3*z_us7\--Ga$]Tj'A,xKrp,2${u>lIO7TDznHvqmA{\TRpn
    Wj=X!1\m#Eu>rQr[5{up'~KVDaa27mo,@'*2eTau1In+|[J[Q?Q1GTT,r'v>s+X_#YHI7#o5!SY2
    E-D\*}XTwu27_{.KX}!JvJ7o'>'~53^0DaYsR\GmA7X^p1AV#na!T<!l'-\WjVV{5[5rECu=,]}B
    ITvr$VJkqcJQlo[B!?,H{l;X^xD@^p\p@-I@rwnaIk*QJ=H=u+TT=mGoJR=wT2Q[3a?njr_UlKZn
    2EEB}Q2*}Arjv#/R3GnaaA\a^uTC!}#VH_D^=u?,2vUym*,$z*~jz{Xk_?@u\wx[0YCT\0Rr5npQ
    r+0[ja5Jjzk5{R\D#_KK7zTQnlYU$HnO!riQ<7Vo2-j]+l;K[G#9UAeHZpZEjRiCE@]!1VXpliDk
    vTp~]j2BG,$$iUx]lDoj9\D]xDBo+6BG{{dQO'azwpm72HQpv~[$v@kx!{r]e{*@YHm@X'p0?QUz
    [^j]zjH*H{7<7YC37Kz'X[[5O<l;?Hm2}Dwx]KYRzu*''a]^.vu7]15mRgUn^{:8m]Vz*+Ho\Gn]
    XE+Oe'OsN\OHR2t!BpKD$A*{v#rv)1V\u~>j-mnvQe7Vsv#^DQG-A~B]j,*zXEtq;CH1VDDz}|Z>
    $vDAa>eU}HiAp1+eY!O\a{sIaER'ill@[[KAQJv]21msOB;,}r_de{D3QKOr~\*Y>1\5/v{!@07E
    >VRUUGs\Z7esI]KIumDal$*TI+wa!vTG[IeJQ@Ia>}yWUs!QD[pZD\*M5J1sl>U^,Wx+$Yo;]w*r
    G?,1R@G@u\\T^i-{1K\pOOQGI'iJhHl$!=$2ATIp}jDVSo[7j3qRkam![TT;}l,.l!==^!*@$kpJ
    :17BV$vv3*Or!X>V$3X15n_RT!axT[CX}"x25e-sZ[a}$^lGUZme{*+aKY%$Tn=oJX_62ww[!]Aj
    )KslQCsx=aa*E[pJYnl,sUTnlo$!ptQS],xKjG7\8Ii$1_?J?SX\DC_Xp~i'j;l$[WO>YX,^smvj
    J7GrJ\sm'Olv}A-Qis-pns=Qnl1<lUa[52<vO-0Es\Ex;ZJ'oxU7Wj,?>Q<[H-vxpVV@C,zulAB\
    I[$r>;z|[>pC=Y>*{v~k2BkeB]!r7{[<~E@m<eDG61l!k3=X$Wsik7}$OOeDuVo>uL{IOU}CVj$(
    >I;THT<,]AQrX+B~zY5k5x!vorH>:x2A[r>z?^nRr2wsYTCm11JTKEiJWYBe^E$n+:b]r<}=.$Ow
    DwQz#luZ;G3H++'J]QwH7fK5uuw$^Tp@;kjD>@+UQ;/l!on]AoHvXv{D#7,2Bnwz[s}JO'VYJjj,
    ]T@>1TZs{IAus@Os?}jmU>e*o<UD!7uUaX;\${H/as;IyZ>uH3{sw%2r~ZusBn~<ArY,ZBve}^>}
    -uyx_rxB;XI#]DB\R}2$;Kl!]GUj3{B8mwj2@j]noZ,51_ZEse5oB@Y@?X]@oYnBzj}u7lTX&l!j
    A{Q{WgBBp2Z7c#IA'kE=K<,aaBsw3U733ZH-[?V!Q1?VX~IH'a}IEr@E-+n_*UsX'{Im*sV5XeRW
    m5W4?V%hJVWK,U<DE{]A<h.[C-Tiej]Ew$+,kOk9$]I#_sA^eC;pUC{V$Qw>n{pYzCYo]zml%UEv
    \lJ3I^Xpo1jsvT}k=oDI5J,*ueJjpHC-opC]oF\#<Vn+5GIm=?eiswJYWln>J-jwsCMT+3wnwp?+
    s;=ACVw?];G]leou*XEFoX>zL{7]rA>R^>n]HV*v1oe?3q-YD2^K_<ZvG2zU{QhXH}T5'V$[olap
    A~<;Y+THn5Hnv?Bme>YGXQ}ZCZWh,-xoa^R\E!>EKOa_^O+{6zEiEI$a~r<ukz]mU,-_<bE$Z$(H
    H,>+_k^p}XaL*rA=1+^UC}*snD@~RC2jLGQx3!E<$K}BeZIH$v?a571[{+'AUU_n]$wZar7;^#]z
    B\Blnz-eUC[[l!{^s3Yk-n.WA{J7kZej4_A2O3UI$oXe,#rQR_5R}aw@-kGZ7!O!I,uw~}KB{@I{
    !rS#\]XzKew;exGrpVpvU[vUTaJ[z_x9pe!j[Ja+=un^eC>ZQ^YHRup<lXWav3eo1P[EkujAJw!n
    v~PO_Caio1p)VO2r8sT{'z7U#2'THEanuopB@eIBBWDzv|@T{@,WAkM[uTsGC~,pe\*:LIYi$*W=
    EWY~u
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#TDnC3pV[ElqnwUJxOKa,eEIYzQ'_o5=}#-YoF"!sKam$zOD\W7Z_p[RZT1us_BU=;aA'#?B
    Bl#^2$+>YT}aap<+1$'Q,AmOoXA31,['>Kj^iY\|_j-RJ+z[lzDoM{vH#&>wCsKhGK*1_}G[-{G}
    hvtIs#$*3s]DAjE>1VXWYWux}7k3HV=hK7a1%}L3,Kx9^B<3IZe_Z[KOEwZXhusBptcazu?CkZ'[
    U+<r3R,{xnGzn{W]_!roB#z}W2_Y>K;5}xx,XR}?x{-Tp<'-{AGRQavMoW2pV{*@QD$2*jDvNJsZ
    lj_Z_}Z=Gz\V]FCKDWWs<1^*2{];O+cmU[lKSE=*pHe?}T=z!fI@Uz-w1TE\weO<or[C#owr,E>'
    Gk}su5YG]50wD#s<jZr|}Y@1}#T[1m{+r7X@R[?HzW3[{=z2]2+;eG?U_v]>B#<k=vpi7Tl_l?l~
    |mRiY*O>1Bkzz^WA[;YRZsU*jTTpEu1#<s{z}JT[lzI7{&}~T=n'5{sVAZuB?[G7IJY5o7'\'Vve
    rxYWs58!C]Hr*i[vQ<T$BY!Top@z7!IOA\DR,UZS#7!l2GkHxImmj;EW5W3HKXG*a=nUC1n*C2oU
    *@~xytEr^$'}DY~HA}T=2$z#AUeev31uRDW[';}<Ox+=W9Qpkon\^21-57e2Z=cJ}Yl]2!nKAzO7
    ;lO1$u>,Xn'nTJ[a^HueRe{E_Os''nGzK,AREKnEz,;zk1x1iDTK<5v?A3~KrCG^^C\J_sU#l#R,
    JR7llO\{lK]n,in,7RU'WJZQ>E72X\W+\@{{THTu[Z;cGlT@C1$53T$~j?mU{p*pmRz'Wap5EK$@
    }vG<q*-l#]$RU!>KOAraO2X*mbT++AgKr,H/S3aoD1e]TasE=w5ozO>n^#I#$?nX-QA'A@-{@#om
    pV{v-H1>op#A@V*{-9W]ls#^!U21_Uv?GA{+zTp;3l?GWa4a\<G}'uv^zr_x3QuavT^k[uj^IGAC
    5o{^xaI0T>uYx"<'EA)7\s2V}_'\7QJ5'vXr?H$]^wr}DIDU<QGE<akQkm-7kYRQmGQNEG_J9VAI
    ;${ls}Eke'Oj{>E,<*KVRWjV=2n*<ZAX!g^w+J'jBsw]o2KGz7z7O<2Q?_?=?zwjsaBDHDIJ-_=e
    jv)U$!]kU^^i7*u_1!~l2Xl|}m!xvI73;$i'#vu$)ww{!DRxC7Oi[d]W*[Z>wg^@<z*,lT=5-V~1
    B*>=J=F*o=m?rpZlTK5ZIvi[C'a~azTXXJ+]k6fVQK_x*}]_1na\<7W&!a_3}}e1Y3V#}2@H?C#v
    uVrJVm@X9IO'nC,K5q3a}H[RYn#vBZis~^TOa$$T_{2>{Z]F1Aro>ER*!^m=wpBk,w;Y=\YEp6!j
    u5]AZr!''as?=;@-7zK}j1JUQBe5$CY$~^{<GKp!ZjUX_j\v-~S---{eEk^%Bi<]vnBGKYiJ57;$
    u<>k?wmvps!]FKl7A}Ym,==r,RXG^ZClIG\*zC>xViBk!+er#>va@az]pv<2Ro]lp-wT#kQv5}?u
    jQ2'pB#IY-]uEp>WzY-5V,^k=l7sT,_2UHj=e1kDpB[luu-<Y7mZZ,Tj,IkeiDa'J-5Be[}TH[Gl
    ABaHeD7YVc,YE^ioUH>j!5k+uWAxB?RQaeY[TV'\+sG'!R@vK<&=OkrCiY~h_G'G+TIH^KQQ?^eG
    rC^pB5<V$m][hq'\XRd,'!Ep_+[Q$~!OxGuzi*5fHGZW*5YT=EVIzx>[@Yv;o}RY!aDHZQ}?0_3o
    uT]T@IRsXehw_[?J><Di]Zx~*^7kY;uel<{W'<Wu_Y7l5I,DZ=!Rs\l*EnQG~z?m<xsmn}]vU@,5
    sZ<YA^svs]nnl>D!^!_$pD](Vp:X7-z7e#H9JO7O:Rjkoly'zxaTB2]G-IAfeK\-\W1!B!*@o=~I
    PlA$l:sFxjB+z<+rZAEXmX]R\a!\>v;KeV[RBCDE5B,a&np*=woK<3=Z[aemGv<+Zd'Tw+TCnmm\
    kXtB;Cm2C,^,7uZ0p?o7rV@X5WBnAnZ}BmRnoG>}E]I<-U+_Iu23Y}*!;Bn~BC_*?7}KBroOV>RI
    r!CsGl-EiwCR}I*!YuzIlOU'^$sCnYr@Y7!zI$2ebv~E_s?=Ud*@H#]"QlRBC-X]mX_1~YXJpTxi
    _7n7C!K3R3=*CA>T'5z>u'>v1{~OGHCI/vwBKI$[{}v>~l_JY2AQW}uH*1~poUeYC2p*<}osamBZ
    15kE!3UHG)TeD>]+_K+Y]G7DnIC;Rk_G=!W'+u15kzHHDQn]v1dEvX<R^zxz]A<~=ZY+ju')5Bu;
    u>lXp_JxJsA>Io+WI^{w#pjU!7?W&WrEsD~~K=$3+;<3}xmCV5GH^YW1[sAOkUj'3p,_Dl@mxA^#
    -Wzax]sn!ICOYQQ]5l~YZTTV^nl5'{H>*pE-GQkAClv_-<rH[^'wJu51m,JDXU-zQH+\$aG\Gw_^
    [9JC7]GxQV\\KsxaHTI[nRmUnB1mwIBDknVO1'SlxD!}s3mr*-]5Z+G2n_ZV=wrQvIjD2]B^@@[_
    =G;wQkrg~GwUhLr~2;VBJKHji>G-BBIrlR9-evjjY>E;1Z!~]-D1=A!)u{3m[DpY,}IC\~m@D<v\
    ^~+p4^<wAoJj;qz2EHGKWTGaY~!7ZY<\E?JDZ]}6siJo>1KwgLPspm_VmG<o3[5QT$Cm[_{Kr\;$
    EV^@}^r_XOiIk{@x$>_73O_{&{Q\pK'o*yQHY=nEij2-3#CDABnO#<V@xrr=GIUa'$?,3lo<W^~E
    uAj-C]OCkD4@H!,mYJJm*~-vAxW_BY7kRm<*C<!%|vx7{;G}V#-o^{>2!C5<J~ln5=ZGT3w'mP]N
    >HXu7K>2^O{CtH>{<eW{{**ek$H'~dgWBmCG<a}Dz_Bk}D#$uXWVmx[,Op>HU-HC'zp=TE"CHZn-
    +C2
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#Ix+]'E5,d2aes}<{#S7le<zuJ,sQU#Y"[:I]k!,>,ivlk]7$'+wnK[N!B#wAG-@<'?2!$;J
    yA7#H#Ull!r#~$!RVN^,]Eemp[KwJUz^;}MJ'+H1vH50xzaR!{H2H_zo<{O^0[;ouXr}x}!-zTS,
    +Q\y>>WaC0]Jr=rv3<N2C@[3(*@K>t1_\eY7is2YI1#5iE3+!u!{=7$B*QO=Q>si\]O=@*2]THuD
    @Oh?-'Eo=3Ec>=$]L~j\u[7I#9Jsr\VIXRO1DarWz7_o>;}JrrVz]'oGl;;5}nR\AkG~[*Ao,G=x
    *xNYImu~*=!RZz3$~pZezv_Pf6\Y2rUaA}CT9!Yi\!RIuQQev;=}i$za7msG#iopshn_k[PmBBO-
    1j>kav')73z,5Trn\@T,3DY[$VuX2R1vK<4}IW3!*uC&zzl@t.kERX<\TJ^o{WCBs<@zE@!T\2Xj
    7TeTw7l\u'us\ln1{B3op^Y.UlOz[15x617vaLNJsWx2+{u$AHXVlA,Zw*$7wI773Gne\Dv[z-2l
    YG$*$oTpZ$+dI+<[F[um\i+Xp{I3!vgZU>UOxK2.PE7,Jz]E=R<,iH_7HRraC2$QH!EX-7>2s}D-
    9)Q_,IHGnW1U5Ut,*XugBzB@E*]eir#79w>W,RGiVg/(Orej<TYaZO-,xYkBvi^+Tor?:rF#r?*d
    3lA_HX}$$'xoC~Zm-vx[YBKo'HV<,3KT_!Q-!nK3XN7TY*ya+Kaj\3Z&D#AGUaoRY3Bj<VQ{=2AT
    avvrwO[<tH$wep+VAv2xKYv<X[UU7EzH$#wGI[DTVYO?-}Z5;1Gr<-Uo22v<*K+j7E5mxj+mOalm
    v}CKkQ?<;o@<E{[sW'~7{-_7lkT<?7,Ax=[ou;<}2Gm-ksj@ZREe],?HW_*G1sa$kuE$[NIoTz$~
    @Z{jpzvnY@V=l_$aoV5mIH,(ps>s$Hv5*iXxATT_/3-o[xpCT\zs-X7+WKV+[FEaK{!'+EusXo5R
    {2Nio1[rnH{~[BD~HZep;pIO,Z<n^Y37lE1\QCXAaB2l1Z}2[VCpv{,?o,Db@Q#s~8^{s#:*Ds!z
    3lp.vBj-_a=i~\V*2&*X,7kXrOE>Eo=T!<}D'Yx)oB=W1aJ+l;\$,[p?5cp^^rUO7~E{}$1;73oA
    T$|!1!sG3KIT$pD@<l7B>_W<s-mBVwZOaZ=I+\k[am7EY]7,$Rs-^eW.|Y@j}$Ye{UVIp;=+HMQj
    T[{{w2re<{OT++DGB^*}zm72Ru}T1a53(KDRm^KH]j$lQ+TrEtOV+DAEzup[E\o!JHPCJ{CT=mr\
    C*#&jW~<H$}w{>KkCej,eEmsnqGl-TowWD3l*^p${51AU[KI*]W*mrA'p1+a\pV~UHh,WJJ<>v=8
    7;7Vo*?\i}1pV%?jk[_U,[CxJu>*_!xo{[R+>EZeR7lQju#]K{jOG#{+RG^o!T{_rR5^w~+OHbvw
    vV}kC^B!5Q]2AoOxI}71;~3sk=yIarHEGOZ;njGQ>,AX{XJ;'WoImwj27ja5XEsDY*\*Dw_o$?As
    D<lY]Iv@E#IEn-32s3~ZIv]RZnwx@\u$>@IUR=lO+-;v)KG$TQ;WZ$3OVJpY$)oEm*o#UlaXA^-Y
    -!}C#1,RIwRw>pI{\k1_D7EjQn#_^iGOBon'r'Tr7Yh{5YC@jRwKAT{^-,Ea+u~}>ARyX]E!HG?k
    el>O~HpTDDa'3ABJ4ZQn#_xX?+or}Mk}]AN-X^Yz,pZ.@A+j[OC>BoDvgJs>CX=uD}pX{i7Z7Kx-
    IT\'o3{;QKB#kU>vp1.Q7~oe2UmQGUe:-o$*aeu<Y<>TJ[5{<'!}#CmXo5E,.z?IG,^?}xvOTMxv
    ajBR^s\vX7vn~ujzQ@}XD[D-=nujj^kliuCQ=?_BKexJpmooz1*<[;*-<J!YZkDHa~{z{5A_$!G5
    1asx27d[?KszET'zZYkcyn=BmC;JIpDZVAH@^W<@}K9o[j*DXo+#{AuGY\^'*~3A=>{BBAY)C_#n
    H\Y21#ww5DV'^K+Y1pQlo5~^rXxVV[olae#kQQ>!\Xe1|53CYUAu+l}ap7-1AmV>>F$?wu|xY{3$
    }n^CJ,@H5;]2n]Zq7p_Wl{VJ)uC\;n]{l$1^;!_2>=oA1{7#~]e!B2'*wEnll,l=JE^uJ2BnEaG*
    3JonZ#nEkjw]Z^?p<C5]IQeJUY[Am'\YBn}oY$GZ3C<vaGnxre1{\T]15\TJ~YHr{]aaY6HYoC]{
    @W=~zsvuJ@1KZ!_mzHa$$lxsI{m5i'2+Z3Z&p<,rHz$^}@lZ2*C]XCK'Qv=uO{<?6\V]UTD)TwO'
    S5!{#D<enR_{?meU\nox+0zQe5/ljJ;ICW\_zOJz_jCi\@;RY$TCYmRCW!<GpK]r~TZ[Rl'U}[A&
    KAQ'!s<{eHOC@O<[.^n,YeUp2,]EJzM:4k>Ra*vB#noKZfDGm{xVAjnxXUoXa]E_=7-_iBk']}^o
    $^ua@=ow5EQRr*,p]-ql35vxIHoXzs!}HzJ\m~ExY*#[G~X?5BRQ+$<qHs]]7kYT{YD?wj2XrAWB
    I]<DE}CEv?CJmo_er?JBoR{7DvD#Y_W\>nnTW+@Ykz~{q@aCUda1\*HGaw7wp^!w-aEk>#d\^Aoz
    7HmD3O*072*2l*THo~]
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#<vKwY*ZCk_+[1@7r^'x<\[@X__\IOz^,7;Y_Gj"O5lD,,5<CH221]5["E[@okVoi=l{j\1;
    12$<uj-ns~{BBY6+1$'Q,AmOoXA31,['>Kj^iY\|_j-=J+z[V;5s;TGX-pC^1&!'Y=YG?5Dli3;'
    p#{<J=ITmJ/[mls;,z{|lOv!$=O7v3BiF2jYC1tan;}iH>Q}y2Ooz,iX;bw+_5[uZZ5QAGJjiVQC
    }1#Hv^<w!a|i=_$$9#>Eo>snIK}AJ?]Z36UsXx!^lI13a,-S[!'7C'Y{pV=mpxA,W}vH!nuTT]eu
    2RX=QIWl+,R1>TKlJ9[%h7Oie{aTCQ[-,pN^~o-Y~'X%1aJz@vi,l,1*@XIjErHABe;xIo$sQ{H$
    =KCrHEmB-7W_$0j}\wG>noR-UrL#p-#tk{-[7+*-{=b{p3@I+<><voBE>nra]WuZ\#wsJCm[cVx-
    3bA1Y{>riI<Ar,D1{]?Xe^a1oUqB;v~3,{]{Xa-55A?$e-a;XCxCos?zZwj!5@])B~BWU[@!uU2E
    *~vspPI;jpm7[}J]Y[p=\>a>p\swlQi$?ZZXTpX{v<C1wKB-o1_<}</M*N<QHU7]=k%I5;k71HX{
    7sEoE;K7pZULRWj7V,k7eVnY<11[[~Z;r=[R_7XIYR!#B^[oi,*<=aT!#XaD>=#}b{UCX?rQ=2<7
    ^}Io>VO}V?7z2jamvjprQsJm$G32?av-Ue{z$_ozQbq&*7<v]buAz5i+u+VZuD|J_Y]PsoQ~Gn~\
    HwY[dhQm$?~-zKAY!WG-PlewKL^TGKqw,Um}3sB$g(eGE^.)[W<lCTjE7?rWE<R>$2pT5>er^~^{
    |G}ezfv'z$a>>W|asw+7tjOVB_UH{iro_#X^]eK>G1rR*%Y+A*3-_-$la=k]7uf}@+*$}u!,7]2x
    <e2,B[':OBDK&T'@Oj>ICYv[uwX$YgE+Xko\m$}uA?;UDwo^KZ,?<_G+nQiC77FPm1*C15#{C'i>
    em-?l2o~~s?}Q>eTr5_1'<H=^sT+iUQ@!]|>jk{ae?z[?33][R~J}?WoV]D=XD}Sm77+,,Bn2r7u
    v!D$+X*Tm*5jlJR^xseE$sK*FLWEBlXjWe]?R,?U'=\@G{BDK]_RmK@+O$?'B3*Oj\lWaGVTK=;r
    xrwIiD25n*I}1]mji2rTl[RB2s_,71}\'~jXuu,xXWqYwI^KT*}a<_G6I,OGo<=U]#R?;1[DQ!,!
    xE]u1EOu=U\,\~XW*CEWY3G]u'ww!7I^]j[u{7jZL[/38(DAwuos+7~'@Grv!1Dip<Q~>AHClmV'
    ]I5*--{<>D:?VmR[iaplW<CTBv'/=-7o+e7Q_$3<qbVBKxNz!p=^<},_NN^n5T7Kx@}A7R7)~ROE
    Z=a5Zr*'*oa{k_#w}V-}'I\]aV{2k17v'o3Y*2_1r,Y?UDVZ8Cz@1sGH7-OEvmx+n<,Cj'^lEn+u
    oj*-nlVY2PG3_}$UZJj5mHX7EW5i}#x#+XOjTR\$rxe>1UIT,s'_e-O[^Z~YWQK<Eu_9/EYi2v2j
    ,m*sCz_2[R[;$rYTCbE#]{jaEDj=rQ,#{]8[k]D@r]vja7?KD+?znY~VHI1{HT=+sTWYGx3mYZO^
    ,]=C5>-^xK!cmOYT%}CY]JQoxwUnCeQATG]{~+=\IS$OD_&zA2mGuBpxE5V]v!^$?2>7QX3[o[*S
    e/oi3;sUrVi]i}YUAO},'z#jB!B_Y2'OToRCXW-jak{B[uAEjKUYUO:{T^+!VwETHZ@eO_\{D~_G
    K\kR'@BIYkxtOlZ_%]I5HTRY}usi5*Ov_X*RKOxmz+H1rGQ~m*!sE*J{2-HAau<{prYu!GH'1HIj
    ir!~^+\^J}!52#A[[BD{EmXG}6xZT2un=x-s1+YYnBAloi2e<e7=uCal2u$]!;,DXX'E*jCRkoW5
    Or>]a=z={E_?~Jee7'r;2I&f$\a$LmDRr(Z$p@DXo?QpsXVjm,,nZ@'*J'sVnXoDJOv!eOGp=])>
    aInqRm'?{UT~]zw!qr?l\$Y}Qr2wJ-_B2rZ3v8aQWZ_WmmX]{p:YXXn1->sxn}[vYo~T}k'}<*z?
    ]n=5BkG@VBYOHH,Css=<rIw|;BY~Q3Opy=wp=VaRk_iOQ^l,Upo];[k1Xb%]QXX0?e!a^Ga5p]Ee
    N#>,=zOmD!h3=n7j3{>+X{{[2O@i-K1-ovI\[Cu{ADI]vUuoS\<+RxxizSAriT-osIz}uVk&Pall
    =+X{u)rkwKtaQj^XDC-d.[?J-=]\_A>I==$i}2_[TpE\weHQEE}<eJxYVtD1_^f+[G*l+ladRD@1
    rOR^2xo_<(#EX>1eTl1YEocvC}KI2eD9eGx=/zrV,y137HI5]C+a!UsouB#Q1mL~jYBvE'#$'ZWW
    -&Keji}5#k9HX$2Ur?I^k>1FpB#nDp5<(oV;nvWvUe^_rYj;$gew<V,}Q1K]~wV}i7C>$?u=nr<R
    YvW5YnB}^pwx3Q?eTu\WDeZRC\d'+J!zTY$pwDo1EWUaG,!2-I!(y*CjK?*R3-annj1rV<=5@^C?
    ;-arx,u-n+75o+IjVT^x3*lxB$B'X\*XzfsuOAk}Bwk'>U]@wo_j15B{eH!=\BSnjw^5lo]~w@3M
    iE,]O'pBfEn'Re^I!rKGxo-=ILX}W[XETe&5oKZ$$k*D{o@6iewlOHJK{H\r,BE[j+Q@Kr!#@U>X
    2X<5ExiCC?GT2Te+~Erx3Glox@*R5~,n9v31j[RpnpDr@*wQ@Bil+RKr{-oA^';E#R]+?5[U?wE^
    $i]ueICHUvTDW&<,Y3XR;TcsBuv'OT{K\Xln5IBD5[C]?^Hupor=K<}$?uOxeZ\wO]?Oe<WYV-CY
    o]I6B+z2*#zu$knAmCI{rm{OqHVDmvJ>=]+es'mHs_Qis6*;a}Rz]o[@'BMz]=;g;Ho+p#rek}l'
    &WvZ<e$}@^o=z$=;De}x_?7-KTTY*CWe_EXeT*-3'3Hw1I+_{lY=2;^ea;=DB|l'k}HrQG*s{W5>
    *sYQwC~Vepz]I-e*AkO$[$I<nn}h^jj1GCw]crQVvr^W+1<>oa,AvpuC$d&~Uz2Vn;C.ITU]551#
    Z&aw~or]*jijW2*nm3($*nm@7R;!UlkGl1!}!,<oQvJU$'iNTGYpv5+CGX@VMmDi!VUACnr#}(}_
    rYC$}@x^?]*2;]X-1_]'p,o1E-=O^UGXu[7_^G|7xo;Y>@v>[5mn'CQ+=~sa>-'@Q,T5{xUp]JlA
    VHo~{^]K<1nQAZ+zB!zwH2^RD[{aY@,2v'o|#Rrnb=[zT+]UWz*AIYT@+F"kpGi_+s<Q~!U$*xVx
    uO{UHAG7eH>njXEH_m?xjDp=Y<-DeRKR>~xp*ruGuU?'8$7^lwsrK@jT1iY*YRzeU<paU]V5GC}x
    m]\^'kH}e_p+].ma\HIl[UlEk'RYn^C'$z4w}!<XpZ{@pTszi{ns~QQaTDVOkjX${o^iv,Y31u!z
    aAZR5Wm$!Yw!rpE*6C,H2|vI$Ju+uUI1OJt2H-lCn$wiD>77#(O_UV[B3'zw=xYX]U#R+D<YV3a_
    <v5W1B*WRx'vkJC!3@WwKrREHo,+RavZH_>GME\@3Ta\RjpY2<\,Go{mlXp]rj'D*FKO}~+'=3rs
    a^M4@E}xQj7VJpBKAwj3Y'-}xuOB'?37z~B=!nr$=Q1@m$n@k=Co,#-jRwGV2_!{zeRkD32o-jCr
    -1{-^J[5;]Oz1#*=jjG'}aUI^eA!OXvp\13!xQ$Klx[zwO~x0CH<#Y]]K_;X#Y?V7UU{lzJ*YCQ[
    nGmevVaI*I5jI-^TKD@@<omQTQK32$3\XvY[o'zk?[p{_s15-V#^R=xkxsv3Kvn]~:I=w[AXHju7
    <#j7_1reC@Uee#Vw_](^>s3KU53o]usG;u_|JjpaHE!@uws3[K>;YCO5Xp$lSjp5_B>5IzoI-I~w
    C${sWBKU3{1KZ~+xjxZsKUzexmr#KG<15W];HO}n*D>\Z=nm<EeX~z]-+nl1u<r=Ew[?~4ok1aoQ
    DBO1^'TBJ72]\;Q=aT1=jvw=J*C-W{=BU!R;m$OVVW'^;kZj'3]\7$j-e@*r@p_mE\>pCT>$<=,D
    jl}j^zz$J3ZY;xCk}VjR^Aw$E1_T<,^A=vVnQv1X]p121@XvO>E2'\BIvE35-G.s1spKEJ=)?>XU
    TH5pA-K?hd5@vrqYa{@ejUwHG[D~DW$WD{e!+unl>'CeD''X}R=d1w'7U,O@;7VuwQ_QW{*m$=Qu
    >-BOe>I#p2C'+CH^~+@B@7Xa]z1~InKnhEwoB[+5^+a<G7iVO>D5V\}KwQz@K\kX*@QH_AH}sJOW
    TB!p34Qkx-mTvpp[vX~awGf}Y5ADAB'-^VR\-ns4,Q+xC@YiA,+W!eEK*?ORzojx?[j?aO<+D2uI
    ueRav{p>aB<*B,<?IH-2pa<@?B1Rwo?ozV7s-vTK[G^RHz#_^V;zVmwReZW*v~Z$,=!*x5TDDW~W
    *,Hl^~BRB<ZI\<e@ULKzlK@Q;{]kT~RJus_A[#r{Dl4I1lR:1,O]F~R1iV;jO|?[#HlCCYYP/pJv
    nG<]*
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#W<+?{$n+DBinVEG{>U1O_Xlk=,wjC}BwFlm[A=@75jYoE;o3*jonBpeB*7!l~Q?-~[pBT<7
    x;Q+OJ<|OZz%lwJ#*+[[o_n=['CW!Ul$HUl=U7BvVO#$skUZ]R3TJh_p?~E.'H~K1\Vm|8Bi,B'3
    Wop?]H?CAV@]=mnxrnT[xVI5,ZT*;[keZkwsQ'_ri}_UA^S<5^$@G-=}>*sI5k}jB]$+wYK'#sH?
    {T]moVQoV#zoHBH$r}@!5z1G)3z[OBn<JBu*mWTo5R$oO\x#B*]D2F*$HO,,?=^Y]D4aGnZ*G!K1
    _GZY-~;Rnn<I?Br?jrp{XU#/".hQwQA/&WCQ77B'i5[DYBB#xc*ZDE2r$J{,{xOA}_^e^oIZGWVu
    ,rIZx^O$n#BH-B+{2?*?xv]GQ$jCkkZ=XuG]x]oGCwzu1^@xKlsQxw@wYJ}F[}oTulR5vJ{Z&I><
    aBjZ5yRQn3nCG$1!CwvXu}=?m;-nA[YJEJp0jVxiGV,Gow_I'Ez7e#B2xeGV12{,7_BnTe}}'msW
    QuV{V5?ZjAV<(Z'J!D1nAB@HJ7(Gz~jy{wru2]AV->B5V3J*#_s'UU@U[RD}e;=-j_GWEDQ@ioD3
    Y\!-'Xjsr}wYT'vb/^>CmQuaTB<{#~U5~2C<[[jiZUe@!sCv[5!72+IkB;}l@\j5zU*?eE?+{5>p
    ;0DmB<^<1YmRB'HCZ=_K_DFZH{kxr\W;]eu]%l?+5VKAKz!<G,$k-\-a^li@3}3OEvW3~1]I!XQu
    #,aAoQ2CuY$^+Pl+7l[GXwOD\iUrOuRA7JD*QO{oK{D_e!tln{uTv3D!77>)*T!?kTVO@sG[37*-
    oZa{e^}XUeuC<5r1C37j^_e@7T-<GCxik=C!_RG=omOTC_C$}SY@7iYjr>(%!v_~!E!\^uV-$T-~
    R+{\nwej'#JkB,~-5xD~CHG;$GX5+*Rz0<D{['H~AB*BQUp[Je[wr1A3@l#T^=e]?=XlV!_@Q"qY
    //c=z3n!]#\l-<K)drV$o9Ho-Z#*w<ereeDi}kk5e~X]l,}2\ojDZWH'.WxDl?*e?V7pi(THjT#1
    ,Yo\*DDwzGql3=woU77%oa_xs;<TVZVwT7uauUV{>1xu@G$UI-lCF^2vQZaXJ!7zXT<{#X^5a'_A
    Yz^#3'?5kQeIl($m{ohBX4Z{~O#}3^#7;p*>p\fv[2vYprYjriCpDIa5J$*17aJ'1Q@O~np-wTzR
    R*VJ_^C=D+?7Zjjx)xz~mO^1']W{<kYB~=*?E#{jmGH=>BxQW|sAE]m-OG_+>vQr_ZQn~U9*D1uy
    uj<Y$#*_l+@n2oo{o9N@I,1aOR+$D]~07}!T,WjBTE,TE8QUAo3'zsZGxsl<<<I?{$I*7E|,[TY9
    ZlZxu*$O{>s2=!!DAT\Bf~\>v9zKCBH],XnrqJ'ks{nrZu*'!sYZuxRE2kj22I?nmT\@I\<{p\12
    -J-m]}!1k\BGKj57>oO+K}=*Vn5=3*sW=6ORkuX=vCZnAv$W2]Rj3k,GJT>^k,ss[@5xXHk5,'UD
    Jx'W}kIr5;lWnzvW-k'uno2eB7[h}vav=iAmiz7ICUCZkV$][sTTl2j;>{>3gwsR;\@@^jBB@^~v
    @eW<,\nAxI>{]=@!RGAs!@73{s?V*[r27'#m#_{{!4!B_~BUwKjgQK[_^2X#H[X3:<>1[Di-Z,em
    1Zo-;^?*+yY]J3~a$klM^{7Df,*1~I}\KDA\OoIRe_B#='OB-OKCw_vOxxw-'N1l!C72vwqz?&{l
    2CkImoiwBm*][H(K$}ii^2x=3n+lJQl]^{K7$rUD2uVIJ]eHT\V'QXC}n*A3E3'AaszrYsQ61G,u
    <Gszzk{>pBjjAHH}~+rwI!'>l2]x_jdT]2[%1@_VLo<;'?sa}+aeZ'!Dj!'E->]V{.@H3n|mYs{j
    -!>*RrA>G>p,5+JJA~xPw7+_<{Q'j2CX_$2OQTD\H$>!zQCHOCI<D5ZG"&WQl!lEaX]z^;,^_jo$
    _CVD#DQ=ljzpxHFAnw+1_UUj7mE~ssRnv#\3Y{kIDi<7>WDBpI}Aw$,l_D+$eT<lXoz=*VV1AY^%
    lMalX{:IAO{{suo@5Tw,e+7RG33NfskAo;$}-l__J\bS\Elvr_\_
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!:\<JrGaW$L^^uQI2A]8opu;)*}1-GH_iSoV$["DuOo>RCw)rj*J<[iTgu+~mCkZ?]Jwp=l!s
    -jAnc>YT}aap<+1$'Q,AmOoXA31,['>Kj^iY\|_j-=J+zr7'D]#$GOT$]G=k2}1e1['@1>iC1TVE
    $CDx*{vKEA|;,~\Iw>-.mrQK'vvrS\HXa<$I[>{$2o<{O3LtKBG$n[Bl{a7>[pwmUHBi{<CEX94D
    }rZ^*\}eBzDSW'G1K5W$Q},r^p}$&*n\;rzW7wTVlAAl+{}AeA1kBCiTQ~aA\D\A{jYGkIZ-HGU+
    \3VI@ipEo>};\osUH[egDJx]}'Q<2,~$zQR^$c!QA$<]]pzvmD!5Al?Uelt[I+}uOCu4'~W=raxa
    }\Zx'3uU;olA)x#m*TxZJJO<pQ'#}VV?B^;O&1W[!^#_rYC[DYz+#b3=1YmTZV/2>s=[;^+61G#a
    #wuwVI7?5~Y3!+urOOA,~smRsu^s'lz@:r;EEn$T!,BEr3}}xfCB*JTaY1dDA>2>*mvJr^*l'#ml
    m3r3sJI<Xep$e2xb\;^?}nYUv-dlIB{@<>JiOJ[mz#'qK*b3TV^Z^Akwa[XJCi^GzK^EuW^C/Hlo
    Od'7w[j}HRjv7DDKQEV5zkXO$ppOZE|Sz)Hx[I$'su=],~HAa@ID{Im_^7D~3xJ]t5ZzD!I>=vms
    }9vW_iN,gGz>a6*RACX[Cl[XZk>=l}8ok}mP{=Z!5?d:#R;I3EZ1*!1!{IR2u<AJ_,J]*UElc=_{
    }7KKA50Z&pwX3o>3[R\~eqP?pkJZYbXB2BtWr}ll5k-Ilw}j?*{jY[!Br7[<zv]rTHe$K7wB_*C<
    ^we\ZCa,Y<Z~U;-z}\u_;}U},{{p]EadkQA=$/?rGv3CkUZsG?Yam11nI]Vr@{nQ1Au{1aao,'pQ
    CjQa=iuA=>/$?AIrR7o+YXu3{37xAxO08#D1]B+-m6d.xIi$<$D-C^A]B_]!r!HE~YrKxDk<!5@-
    =^x!~^77w_(,~Y]<o1m\@Ii|kUJ!zn~l{]\X~R]VlmoD7]EXQ@sjZOza]-vuCB#aK-l^ie2-<}<O
    ~$v-uBEKs=kVve5+O{maN,;XoNd!B^@73WQ=@@E7~-Vpp\[E*rG#Xs*[}p(>_7,7BX~+YYr-$jKQ
    O}7Bzs!nTBVr=<Q01CoZ^1jBB;^'vnjVlvAWh1T\WPQp>WvR[l#B,@p~a_^OYA-E13*=_~X]KA!l
    eQCpG7o1)7UCD'uBe?<a2GK]koX+rlu'Ez,Be73]7l}]?Rz=n=RXU=(1_Zw*GV@CJ=@1Hv+l3uXB
    IuHN!DusD1'XUYIDS6{X-ZFGpW!,CzW)UVUoC>{#pi@$%^jm=8QlvY=uEZ@}]*I?J-}]IOHEiIV_
    YCo_oH'J\>QY@v~Iip<wa=bnCV+DEIuAH@7X^T<v0]aC<'>T}G7QoOODnzBr~'e_ow8/p~<avvKj
    5E2BExA+sTs$AnY!G#Wv1-,XD^~a7VTXTA7=6sjn?@RIIb}B_jUVX=7'+>.>r${|1?3sI7A{aHr}
    IYTQ<s{~sB!zLawqu7IEORk{$Z1RV+2]eZwTOaXoVxxr5sA?mpvUv1X@@lv$52VZ*k1]U,><BvB@
    'Apmi'Xol!WGkv!KitTTD!1~^nU9b'&k}{~[AUoDB_WZ,U@\OjDDp\B1HowYE{oV^~-_kQE+*H+a
    =DH-13C4QuJ1UEe3'2H[2ajEG3~5C{Y}B>DD2n~a.}@3B&Cw2xW]\^]B@K9iX$_}*}@z7]J7C^[X
    {C'^#Jl_nVCC)=fEpB'T=Z!]EowU->{p#,G>17<}aDi'8x5pz^Q3+7DDpYjQOran]l1>ZZ,mEOxT
    G#-*K^ZG~Ex]BTvv[^^^T;Do'?aQX]7O{ksVl|v]I7hHCneGJ{OI1V$$?HOJEXrfD^>A$BVzgE*9
    8OU}@C-~-[@z;R57slXx5{\HGpv}TeITkWjzAc/_+[*K<arr<5;\1pVR*3QE>X*@[2#/1*E!Uszn
    Q@$uX7[Y/k7pJpi{v\3,QAG^zkxm$sK\$KATlO]-z6mDI'cT]}O,iplwG\k~]\Zl<*pp1{-{>3Qo
    [E{kO\e;-5CE;A<L5WsR$@HUj-^ZJYKl^^@~OHGJOD'3]M;eV~?XQ2C?!+@z5$'V*@,#Ds>pl2rs
    $-D3>Aznm>*W^E#E6V3jHHVJ?E-},>ns$VQ5J;>1v6{+;a^H1i7m_Hzo{<CDs=Y,1_p@XwwX@I>D
    'p}Br}^7G$\i$Bo[E},p!3-[Y\~sleQ+l35k^o?aXKw|K7$x!aTH}iZ$e^iI<\i=K}sIELs+C!tw
    _@z+5G#II1@<erpR;rEx?ER=rm\7,kWwVeHIpj3t1$x1Q#J~c'K=#O\_E[#Vpr|u'?m[JQ#,;!_m
    *v@-x?R"$KxKG{]K}<
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#,+A?C~x\vBI3eA,\5l-R9,BEvjxs,ve^i9eCJ[6w+E[J1pA!I;r3emU>R57AEl}l>W5I$;O
    $Qa;/S#Ull!r#~$!RVN^,]Eemp[KwJUz^;};<VnzxnXXA\JxYipm7#@[mUw,0D;W5r#DxRu$#s@7
    [p*oY2xTz?H'I~jzZv>m;|Vur?IE)a[D2>Xz[BkCE{Eu-I_elZ<17A+0Fx,p!T}$UEDw;]*Eru'l
    p~T{E^'T\?7+T1v[BI~e!bfHAY>b^i$Kfxz7-#NHO-T#w_wH\^^mU'R-}],Y\Y[|K^u2+1##'O_!
    jjs{kXe%eG<Z=m]aIB?3xIs>zm>ka]_5Grk-m+[~{RO7Uj<+A1!I*,>C1x?'=iD*e$uXQ~{Yz_=1
    ]BV>tEG-,Ql_GE2p[E@ve&8{B_px@TY^>[AOdHx;]}mI_"=^KVsr#l!{_@U$GJ,B^-e5a=77j@Hs
    I53DjYiw_ODO##lwQ*VnQ5XEYX*}QY=?=p=]YD'Ro*\lOUTrHIwr2?^GRa3we_[?o+=~\s5YpT!T
    D]cek\^5l,ikhwIrRiYw}\wu_*$wWY~GDe5T#VlaWEouBrY@s]^pnrB=O>ws>jnGGXEY,VU]x~{J
    !ZTG~-UYaTTY<=s1jz!;>-XXrs5oQPBWA^#}#T'wJ[3}_~lHUE=5kr}isnmA^@
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#X+xsenKJ^BREl;1>i-o~=lwWj1k[CZBw}m{jUr?a<T;r2}l?e=mWiAe3*NyOOm$r-$my?oH
    E>5zT<'k$_rPlwJ#*+[[o_n=['CW!Ul$HUlIH-BA=O#QET}7['ITC'isz4GD-n#]X]+Dz}u[2u[%
    1xI7G{oK9KhRjW2@R+2W\p2'r2k$w=RHV=io<Q{\Vju2GfBWa?~UmElQR}>^~Q*+ETIZ1roD\?YR
    *nEBAO1aZ-~AzH=@>_Hlrx?-E\faXxjlxQu_jGwr?w;E{'Y7wQI+{5BR^2}pj*Raj-Ge/W]'VY*a
    A|F'pT7^XEZvRX{,,I25aK^H]CeHo{l+A*$W<\T#O^1<wT=/Ua-B=Zm>Ial{QlX^D1<mwv$+^lX+
    lp2OXj+A@_AWV;Az$=T-m_<=B~'#QD7OAIj<:>QrQ#>R{is=u>v!UQU~JOvO18I?!sk=7_u]V^#^
    zv@<T;\ev@oZHs*rTQEU+j1^n'nRUB3RaW+QxR*+A~&k>_r]3pRCZ\-tEVj,RwnB==Ckt_l2oG[#
    BJr!T?$<m=aRKr+eau'To:AG5$*:0_sB,g<rQ.5$Y[]ATW'-luj[{\_kVuCQrp37opppxRAX17]j
    ]pQQ'Eu[~30'<{GkTWCZrT<BAU>Noc]zZ^=+zpliVZUo!m2<n,3-un[\J!$Y;z,4QsXzsK-s>es{
    rDu$lAUI<T'-^}Do<5z=]O@;~_@HIW2pKvEU^5e$;XzA*aa;;'\z#evX1J=oKUBn#j;?l!3>1V2G
    J*7QIC2],-!OiYi>Z*Bk0lW$Y6kH<TYnX]x#XD(#A'5]R+QHR'OR]usZ,IK{TVUnU@ns32-ITT?l
    KYlVaxv>UKxpC\n^D1Hvx7pT+lmQH$K]E{TCOv@p\p>&?]m\3*T#Y?aAW-J+S_=-a*?rpx+'\7IK
    \#eHK>O_aeZJXR~aUXR};?}^>Y\uX!=veu_xB1_VX,5_;z[m_J>^;}X$m'-5{T,;,}Xpi81-wsFd
    2$~1x3u{K{_HO1a;oK{,IZRJ\il<!{n@#xmI$!Hzj^[A:>,wk7\??prpk1Y?e~_ap>-5B2IH3Wn5
    Dsl#knETDDuwIk=}KGwmmDUmz+'kw{}D?*!CVelaK<]=u,{pT#V^J$u{YI?w$w,I>e~@R:wHXX=+
    +=#}*DGr,*Y5Jw~{R^G<E[8XO!}"!Iu{z~UVQ2W_[B\}Du1sX\5uxJKT#D[EJ{rYjC]?>*Y+PB:#
    ]?s.^^I<ajl>N3$2Zq@Dk;^>HBBWEz/$n'2]$?J7e'$'\A3mo#,^i{$Lr,2?-wU]&wv};1U{]}v2
    CHs57<G+?@oE!G$k^RBxo*@z*5ROo12+wyH<}z#YXURQ=]}33V5xDxxsmW/vE~@ADG>cB+B*J'Dz
    lIU@onU!#^5!lRHY}_iH3*$Z'#]uOT[]ZwX#IOD'YE,CseVl<Dn}[DA^?nD?;1ARR~{pW-vsJEHr
    !Cuz^3mxO^jpm+n*XCZu$^kx_W+<~}Wa73Y;$Xowg)T-op:BpC\vrJ1mU{zev2o+G^QAG=U'Rwo1
    -3lCi32^-]rO$;CGBGpYm>eluV{=v#;^u2wGe{+Bw+!{<A]uownlH+G0\\^K}e1*zBGss@rrWa2@
    !r-;V5v+OGE+|^x53Is[}ekp1po{D^,j>_JD^eW\k\oZY\^{,jHlJ=[-\[,KvjL$iD#_o-@?IA@m
    U]sfjI<'U\_-r$2JnQnuBVX^C;$!5,_a;oQesamGHX{uL@{=1['A;W7?]X1ApHRVB#C<25lm1}q_
    EB1E+ejJr=-/+=#lwTl}Jx#[q7o1re<jR".$[B=p$][_K+}YnQ*Y$[#\Z}2[;QG$x1?D8+_OimUl
    i+I#!@p;7(=dCDiDKzHC^NCR}wu*{!junTI&uQ*=B6~*Arz>DY\Z*JN#C}RT^=YCaaWW^k@xmp_z
    ;7k'JWsv!VER:E&>=>G^2T<(9:I>O{{zm]ujXv1A]W8DAXnH^{=zQe2,rG5B5[vAO$WE3$GX7W7I
    ;VwKjn>2E=o\0\};s;Ap=vhd$sl2l=m=}_{n1$pzX$3'o,T;t(DO[]F2]!WsZ1ZH+{QBr5zQ~\3[
    ;<JzX$Tmz+B!_A1nz@'[us!>G@k5DEnJazDur2xQ~r[L8*|~CvB1D<_\=T}s=#Vup[mRzx~C'j1)
    _\Zm}2^a*\}Bu\[D$<*TC=[IIf}mHUG_k-#rusGG^RXC@j$Kp5p3U2D_nE5IHJT\JDj^1l^jax&[
    ]Drp^oEB!P>Qw}xBmnpAGY7mBZn5pn\Q<Kwv}raoixpn1oZ7\O5w^QR[5[K(2rn,o5kz^|YDD~kC
    V<G\!{pK-Q]OT#mCo}}QOE;l)\EEluAa'MKEu<O<J}Qx>o1JeOuB7CHTGQ$7H$$\-vBK}KEwo5mH
    <=_^]7!*;U#_zJ]{;JGwpaEv\2lI?1+vh$W~js2_e}XYY<HTYYl_7;l&ymB-*5RCu3$A;+7K@2Bw
    AnU(o~v1JeC?NG*$uB{*H{aY>J=H@Yv]G{5$sM[;~@[-Q;j^}C5vUs<D$rQEI1;7kpzIw@2+;^=p
    V2#r{3J<a^F}1mZ<GCQnww+?VmkVzu$r7{$kR+I+55Y]sG$UarH:R'OiAq;>j*C!a'IeaH[}p;3U
    ,A*_i[}kI>L>EiV5s3J3UCrR^>jBu\$1!<CKeE;$;xK[,w=<r7I4^D-T?G+ZpB3vh1vkpDwlHvlv
    H1{H3XGzV5UZa;r?EiD[WcT7$'<Da\GEDV;RE2J<rW,'[3a7v+OnpXzX!s27\3p;pYqI?uWcI\\k
    Y<~'\'<3DsBBYX<#Uw>~+AQ2DnBJUOIes$oA,7O$kn[vIg}\I_BY7sUpD^$|z@szCx$#Wj{D'ma;
    C>BkAOv;Ha^I,#Z23OzE-+BQe5}3~A}Q1W]aYxo[/mQI@aCTjABIwgKr}WpB\hV@$=J5^>lTw{p.
    I2j+;eZHE#Bn*CQma5uKG2{O~a^ZBC*#~a$7,Dsij1VR1D'nnHw1O]5rZD>D),KJXVnv\o+IA~v=
    RT'T=\#7#$3[kn<ooc}w[UcAn5B2CZGn<}=*?]{,*eW,}Z{e~,<p}m]=+lvGs';C'!@]nXD@D-[j
    TA[X_>lMGu^1-I^Zd~{X\1w-UeaJ~J7\H-jx]B~~k2BKXrTlE\ixRoTQ{uv[o"XD,2xi>KO_+B&\
    k^WIz{5Tp1nBXo}B2AC-$R*xvZ3>TO[eXl\JvXG=~]vunla2[K_Uxexne5ay]~\$>^[eo2Kzwn,o
    ;^kVhE=j'^p3ml#p!'z$3xHA2GHV=;>UE=o,'O^,'ARw+ROe#$]ox$oR2?YHo*Hu7wx-,zB@[;Rw
    mO<Qxjz^YKz\vG#vEvH!#3[]@<Hs@:jXa\\U~_EGjw;1ov=uEOC^~Q_uXU\Jv'=\mv3,@QnEvQHV
    IaqxC$2un$T3{Y!QHE@D_1H!oTnvpkRuDQI=*XExB~j"-77mVGRC)r-^=,-xo]\-RAGXDwDQ11p=
    #z217#xxK*--B)^>VXEYxD=W=@-B2CCk=pI[AHEGa7kOkD'T->),5_Ey%jDv;pHzxp~]<Ox~',>s
    xtWBBJ@w^ZA{^R$Y{H$D<T1vQD|G3*E;AmZ6^{nA@^k~o_73d=m2x$J^A'j712=*EnY$ox#HV,?o
    $IieWGHJwzVpo=CU**}1Q(d2VVkIK$HUwv~kO^>}!;=J+r}5G=$Tr<xZB$^ZnAr"]'{5ECB13(o7
    v;2A'3*,*70ar*pGZ3@lo-2_ICs]w!nGi;J9+TI]PGS3CE3YABm0,YOK^?>1On7l7k=X3lVB#VEm
    R2JI-7pG!O2[]zT*$[3+BK$\ioeVpAE\xX~*&e?swUUKXP]{s1i-+>j,\E+T2GlGKo2*a\;1mnV>
    UaB#B@1ipp2E+=PU+{m*i,^$-Kn>+uY8EuJ'^OA2{=IW9z$I<ssRsz#GjvV3ofD^TmR#A2pv,Izm
    Ts\]]iwTp$v,pW1eGU~5KzOJ^e;v;3?YI?nRp2Y1R7[ivwma;7Uvz2e#=~p$_sY\^=^][;}KGivr
    ;p&iE]z-Tl,_eKD[HjRk5;GZ1v{_~J7#VV2UA@p/Xao*7zv=BCIIms<pGp@{*{@JOAm>{$YvTv)G
    _+o}}I1a-GuD'xniD_i?<owa_H@;Gj\+}YEOJx\V*T'HlV2UTErq}jeQXVTj/6YT\kM\[mQIe{m@
    O6',x2[{JvE?!jpaRwmC'p]i>xrv^px#ouJUWTG?>lB@@lG,~-l>\Jf$WE->*K73<*+~'\7]*JIH
    DEEu\n]OJEo*Ks[=I7#q0ACV<Ax[sIKW~^RWpt}so~C#lKx3pn%svEvwl<_?ll#:'TTZ?p]}x-wA
    Qu@u^OoG1p-Tj}u{I#$Dn*,-<H!{~wZIvmln]$CDZADjYHwKx1EvlzEO2a^DzQma>xxKq'@X=m7!
    G<+TGDU3oxiVQTr1?7n>U12!Kl{3{W=XKl<[xTAn?cv}T2xpYK#$a23h4Ux*=:oi}U)DOw*ls{=r
    =^Ga_iW{5*>owwI]1l'T'2jXvGC7}}RHBs5w]]U*C1#&)UaUOJpE_q@HE1xDp>-B5W4;\!keZr~_
    >Uv#EeR'5A3Ikp*]-_[GDp,]Xs<*@;UuYxVECI[[{$<LeETODEzx^!2e+1a<Kl1K1OiW6W*m\4G<
    +uIl3AOT7=zQ-#sXm{*>a<YS753~O#V!H]T>-,XKY$E{((J<slBsm]?rGXIHukWQo_=}*W-AG}\R
    7#8u]7-|wA$$\^]!JHDW@72RBi,*vW^E=!Ev*AEIyoUQ$e#1nV=<TG=;<YTj_^dR03-ali<^De;C
    ?9s^ohB[ET*Au7v}!D_DD-'^_<-pW-W<Q__1~CxmA+o_w=mT=*P.*5[zJeiY#p\aJ'WX1>V>x8]E
    Ejo+Q5pDeQmjTmZ{HnJ]<I:uU\a9k[=ww*KG_<msI]lHUCaOK$eBMZr\T}]H?{DiTV5_w*]Yj}>m
    UR[,K[]K{C,@[-UVx+DA~<Tmz:ojYGQTXaVXjHv?-vR12-.{sjU*HUUV,V!v]V$5TC3QEVI=UCp=
    ^jlVU,@$BpRw1IY\i1RzpnvBUjTeA@xjanjRTI]WOUB;o$G>v\@zlD3wEE^j-G}u1eu-OGJoAKVz
    u=ko?lWQmuxnn>!eC3{l0ZB+~7;oosr>@K\G]!5vsIjHR$CI~$[OeeL-+-eO\=~B2Y]S~O!;0m>]
    $f$Y**B4_To7GJD#;zT^=l\<&]1>T.OVDGr!=?zIjOvVIR#U+^=['VEeHBB>~!U_BA\knw-^Ea3n
    -pRa<n}!jZBCEJk+~{W'e$EzBTY<D-275#v++p.*<Ynz}m!GusYfp\?wE=o+A[v2=jjQ[u2<I'3v
    gAjn39^T>W$DRnVDw+pZnE2}zDexn3T^Y*WoZUI$*[,A$zV^lY*wx3>ee[T|~YBuZ[5BZTrukA>l
    -wvvK]a,6.eWW$x*{_,ianWQ^[TELiUXk%~Ga@Oe}C#^z3l@23b653z-%BtCAoaBGa?_m2p?YxO9
    {q6~5?m*a*wn7DQ({{UZ>Gm2j2_J=TH'_{-KIwvY,]=32[o!4TRT][@_Bp<YHzevU+V#Uo]1BztZ
    <AjjZ=VVT;<s[nT;XBrEma$E-j+rK5[?CTOs,1Un<_BDUz\'U_C5RW!B<DaOOA_{C*~LsvBKUsIY
    ;{B2va,j^\u{^7AwV>ZYziH^SUa_iw7[+@H\$I$o~RU7JY@sWVi;1c'^Dw\n-,/k1XHs\[12,uER
    *vQ[T=w=1ne{DI{qk>rG12{;,^[?G}+]|Q_I*q}{GK_[$Wp![^@v,KmYT^'3vA(Bj*5pu3kqYRr>
    -_o>~Yj#x?I}Mn}HRT7_@H<-wX<+Iwp_2J+eTooYp[;+!lT<XU+E^A\'!E21ovB>u=eA?'oBw=-H
    +*nu>3ICu3+T<sZ+21GXUrsAvOQ_xoUoV%!lwl]BQXW+5#osUIBIH1o-^$xaZ+mr#su<Q,PqUI,K
    xraWxT5]AriTm}]k#XTmC3p+x32eLYG!#CX{+2+anhg,&;aJT$Ijl*v=2RHEGS7Bp>+'e+nX2jl#
    ;35$$^jaUCdGI=]7vJ@K(xSpx1k+Ovl+s532^Y'B'_V;j~j$VnXw-'~WIVls'*75vw+mxzvI1Jos
    @X\b-wA\Z\>pB=RsAo#D(O^Bm'<I*xGrTKIH]'+VmPwx5Wj+;sTxAKu+Ho?_1$,RT^Ot>j^<e-O;
    Ge#p{pEk@_Qz*V$iIZ1Ja+-',uD]G'\v9BBE3ne2vEKBDre~z@=Y#C5DG}rIJw<Q?+*T751$OZT7
    ^^D1K\]DU@+j3tPa*XUHCYr@A]Yj_s>Y@oAYzz+/H}aAlYv^EDlXo{a-rVrA'I}K-5XxM~v=_YVo
    a{+l1je+vluj#ve_@?<Y5Zj^v*,T]7*~]3'R_DYoOeUDk2E{'Bv-UlQR[CWu}>'!l7,jxz<xiBZ-
    {MSr3Y#kxDRn\R?1X-Vx#>T!OQs#,=2{p\+/_zj'rmU?$G#n!CF^[2{onY=B~u]_r<pz3e5aO\*u
    pz>X<DTvEZ-QCW@Y$#T>j1oCKOETx;uu^Q5E3vv+}7O'=p5n<+C;1p'_w-;=5oJHwUYuA{G:lUVl
    $i7CvGlYy$j*1^v}-=^;@AE+;eQwVe]5Yoj1Q=s''["_zE<IrTA@H2[D,=m$O{o\Bx@jG^zWokT?
    1XAD7_~5;\r)Y->_w}[lUUAKie[$uoC\\w3ln\!<V*:x~Io-X57QE7BvuIag\?^GC<I+FuHwCL,j
    npvo7Ij7,5u}+]BZVO5sV+^7Vlue$;[-{~V>z^b~+Xrj^<wCji@iT<#lnjoXCnC.RW![VRGDJaGG
    I\,#5TjI,oW7&VEY5k{<=mA'D:C'Z3Ce;=RQ_!)L]]?BpmDpS*V{BpZp7|7WRnH'mjZ>nRv*n_;l
    [K#[<-AsJ>~s>Z?<zno{H?X-RU<GT[125_vr*=]x<UeJO#]!~;>viT5ou@2AwC:}UQ*?=p7o4bia
    uIj$-k[I3sh.*3~'/kX!*O=O]lZp$O$*Vs{z{d{Y@U^aQu~onDl+CeL-s#H<B}!&@_X[IZ*s%+o?
    \~_,Il}\>aHm3DaE!r11$s5Ds$$IXKCuR=]I;N:E=\<1U2Klw_Cg<1TKa^+^T^BjUou$oYX+'J~#
    o@2?~w(3xH>RRV\e1\AOT!E+{rn]m<*tnrCoHwx[LanKxe'x,jX]wJjz[l.>{5A#R,DO^5v2XCKT
    T{D-5<^vU{XBmp\m\=QCEG@x{2>OnI1rlHa@s_@<leiIOE+,2'e[BVUrzE\{5*OC51G;,+p>C@O>
    {]Is;UR1xqC@s^_Cjr!jnoesEw]TR=72oC_zA3W7=[\}#{=XIv{Y#vmY#H]f\KG2G\AGc+-pp>G+
    p3U!vKVwU]_-RZ-I!{ap[\'#C[O[T^Y*+BEX{91Jsv^Sp1okQi7m99#}!ue#vEiU]'55oXQwZCAX
    Y_5KXpo$\De-O,Cv]1#,+ReZZ-I!!RI\R_HsX3AB3U&kei<Q__O=$@wsOXBZ}e@K+o>uYe?y=TXe
    k7DH'lU-.WlTsZ>7,@UVr]+jwI3R]7AZRQKVD5=5K^l,pE;pk3lzlj#HsI<H5^;xE,>++:m[e1o]
    *iR*G=?G@@|n{Q!C)Av[}{Hl*uY;x6<j*rX5#2[7'K;G!w
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#us}IIm1s!X_u+Ox;zIIlYTaYROO,+R]Z};{RuR#UYA<sw}'ViH_TT(Q3<<GD,;^3O<|d1\}
    EkT3#vHARvjk}]irz!w$wIi@DFzx^QI}VCX$sD72[lNW'#Zz,#_{=JUwO$Q'Az~wa*C2]^!*A@~E
    BBQ@+YBzJ'\}TG?Hw!$reUw*7OAi55=+{sY)~Tn2'G+@u,A>DiWzr*=Y2BVp3$)<V~n3B@H}i~E[
    u2?\Q5$@C[A!pXE{+'uGx1^C3uV}j1U[\#xJat^pl=a{jGHx#nYeo][G[@i-'3]]+j:Uw;X=I3uI
    ,j5Hz,asC?xjK2zD2e-UD-eD=<$/-("DI,BMOABH@1ln=;lK1~3I^Q#\B>lx_5lX~I!',>n\<Ooa
    eXA\WT~$wTH~1BOU~s?B]Z,p<Tx^7>u;7nuAUH$T@o;!U*m>kB*j-{BKzVk,O<piRlAJDsAw!pE2
    9,mH]lJ1Z3eVUR1EY5IsEWB]D>wKw@V)<r,Bs2K}iX2XPYwUAk5K#<el\N{_[T~Hl@Y>*B3s+}Oz
    GJ,i5Cx7R+v<l1zU-nRW$j'V[<6HG+W+HXpzr-o_xxlWYk7Era?.7>{jIJu{'r@QBA[Y|Qk]3x_j
    !vN=2DX%KTT}z$A7L*Gj#{Yu^Kv@Dj5$Q'Ou+pv}{p\vApBw{}Ku+Gk}@zk,<DZp;1GeEaYR~!X}
    WTvn5>Do<pQAB71lCYC@CV2Y!TOW}O}[}l1p-+{=BG>U@r,,I)5Z4CaJOOrIG+G3DziQ?ur^7<D]
    j,vUnX$$OS^T>_{De<]_!l,+7@'1,U,~vzE=}l7wDs<^z!'p#mk52w?sT@^\G+-Czv~V328]Y^rI
    p{@2hJj<!1Q]<vkln$OOD@o3]Q+v[V#uC{\H>{7
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#IpG5'Kankn>$TQs<VEmk:\E!,Ewpv,RY[C!=nF"BO=Y>1Uo[-;Ubsbz@X5]\5QjU37Jr}?e
    Bp#^2$+>YT}aap<+1$'Q,AmOoXA31,['>Kj^-1V-]3]_7[{jx+v}7Cmm]nK*H{}jOE1|,?<@bjT@
    J=Z-2}RpQ<O5[[D3<hxAAANh#EV]n-<[[BJD*V+$CuQ]O-aDB}[HwVrk}]Q7$3G@Yw*Y(nSK1u]?
    +-ska!Z}2DEn>pkDC2ZhT7C"xjWe~jH]Gf#XHvF!vBz}Eu{Y#=W*_[l\-Yi,kIZlKaA=:oT{W/!O
    JwNI<2*}Cm=IVI=U[G*^wsVqHDk;ZXpx/5k+XzRAu7?Y;^JlEJX<$^IG#$ulpu^ZWp$>_$-GVl!^
    aFwIl7@GoTQsU<<$UZs>wR>xY#V^H?.%kA}s&CX1EejOX,1-AkQAC?ww746t*,X?UGXIL\w;'fBD
    D\;_z],$,kU]B@s{a_,Aoi3e3jH$EpIi{OrU@-KE]B_+A*2EZ,ov]9eeUrZDnxlmo{L_WR$QHY3B
    iZQx=zDZ^>v8'zxC5pV!#<>;2_^}Y2Q-Azpw\*Q,QI~\RJ+^,ImltKQ_vf&rD+${}!*#N2__^@+~
    C4UQpOaor'}^rCTrX$CI<v^pi{T+rj72Cx72UvBHm,73-WUv=OR_Dox#nH>Ri[#v#o,j{\!Vle#7
    k7zg1[!c
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#7*T@A+l7YZm[<T2<$;^,qu$BU88YjBr7m[+-]i!ViRuOox*wQ^$IXHDpmB*p!x2~sRiI;TH
    {}no-lX2zCC[EfkQ'Be-e]iXa[zx^QI}VCX$sD72[lNW'#Zz,v+-}5UCO$^,*?~~aZvsDylv][I?
    QV[X1Y3XTT{T+{ylII#iD[_}WmnYD#v{_jEd=WZJ}\_zEO$^{siBB,~Z#<>rUr7CKXKsb-}@mXsI
    ?VxiGqevoGTY>r5<WunTD<15U{|f-rm~xv2I<YoDpRo,~<Rk-AW3+R[\AwV2!')=^5G^<QEp<Yer
    ?vK1HQYb^w@;#|X[{om[3kQ-;<]5J$[,RzY)B#[#:DHXov7Lo$=}}$Cn~=7]v}#GrrUU25An1nm!
    \+jK>7V}YOmTK5+G5{VQ;l#D-^OO'U\E_#ol2SOi7Ykn$uB!Z[@noYEH_7bV3[=6xA\]5#I-Xau$
    EG751vuaK{5l4Glal.We2w@Tez1An$m]}uinCu<UR57X_3bOXeG"QDk2$C~@D1zBQCXYAEDYp7Tl
    vKlww}$i~Gn!}HWDx!VJ^Xj>^I2#+E<HX7Az=G;1c2wz;v]{;2C!e?IRGk,YOG5e5m,vX-qw--'0
    taw<V]Xu;lT[Gj#QJHjI1Q$>YmjW<nQKW9^_J?O?3@#_2xM3{XO@*Jo9]1omC{}O+>J25ZmjpXW@
    wACi\[s?HYQEOV#D^lipel[aT[BC^R[z1GzTl?j5Z'?@'IkCmw'X^n0)lvu]~o'2>EDeh)R1\!=$
    ]]>_X<c=\]Ba5{G^TQHKe~$Xw=@G3WGAxE7V81;JzTOG2xOJ]R1z@AX$~*>ralrZ1u\zJ3=RJBrR
    !DJK?T1xT\Z3mx+$#nAaJH>uVBZT+R#=JPsHw\7le=z=z*$C+OeH+oYs>~\2a^7A~\#HE?n_u>$r
    p+c<Ik@7@xU@<lDk}jw\?lG$n~Dna\Cql-VD[KTB1e<x=ADD>AcT$DGYH_m-n<>~eR*s3^C@'_*p
    s$BBY<AVr<K:j*?p|r!w~[;w2EHB-B;Zo$l2=EiGT15{'=r,uazsuJw{{\Z1kZIY-$WZIn5z]Z]W
    1MrV=e<1j;2r!!KaU!d'\$Y$=pA7DBs"I&#rn33TXET-61p2X=HpT-DE!Gi;*zeC@wERaUT330f7
    _$Il_EKXS@=o=,sj#CuZY=zm'[+x?v*J=Ywl~$]mpa'V[QD!XID-rAlkojp<*(oGm[}G_m^Q!u9}
    H7J[BK'GpAuvB^5l#^@p-2^R*a\<RpVflmrxOxDmKD@YJ>C7l$r_H_QA;n-O+n23[5?$QOVxAR3O
    }p{#<}x7^VX^p*iZovUDyHawQu(u7HZKICl}?Cj]^}CLbX*!nQnG-~Y5;TQHv?HJw?O-KR{WV=K_
    TeOKsAVQeGDT'QVU@=Dl]',JR''HzAr,@2RXroz~7k.C<AA@AwesE_\9RpY^l9<rHz\Q!zx2]Z!D
    YKGQ3Y<$X=;jp$DsWn$Rl5'{w?FnH[=BK~H$pnsH\=Cw1\+^kaJiUBwanuj%rQXwmlRzO0>=EpEx
    l!p9]HvD~VjO'm<Q}V?W:&<vIx^XKor~Qi.4v'><q@DzHO<j~1-Iw^A1OR]$!_)C;v^Qz71z}mOb
    IW-?aQ{=^jkp#HxioA~=$mEe$anp7U{_[nIwX17As>sp=[=k0$j_{[lQ~E[YGAXa?E3AwTO~,eA2
    GH5?jVIUO$YreI*anH=_#mDTaBYak1!Xx|C$]OrlJGa,u-KYX,K]]?7}uUhy\*kV=,[v$Z*Gq%Jo
    s;r;+o!w<W?^\;pv.hRlIA}Co7BT,mfmSUo5[UVc>s++x3>{>Tm~V#z@B_r1q$p!vJo>}]5\D<v\
    =zQp_>,-a[;_CzJ]x-$Yx/]]uKAC<X.fI_oBVj?^?ezvDluoH[J[~w$3\[H=\<YC%z%q}^wx1a5X
    xm7?YvR1UBA#zCU>$#\kwRmIA_?''~rjmOjpa^m>1OVsZj=ANe[_IU7OJ;R_ib7H]v,JWY]7{R9D
    Uae7\Row'[}B!@$eis3ao=2xI[Xk<~Y\>KkRzrsInE#s*}xDRXTp_!niz]^O>~rnY[AXsw^uw][a
    r7I#DkERJJV?1UTXop_A_;ZI}W3nEH=KDU+RuH?rBB\}>^]Rl1$R'C?u<zE1ITIxI2'?\<KRs*\r
    XHIYmJ3wnTU}}>rYCYv,!QI^1eEYQ_'7H[VK5<G1pKH^#A;j{DCRB2n-1H^!nY}m*?IvzVnIsw]$
    iv1H-VUeBvC"->Gu,,+B]w\J5V^'3EmDA'U>+B+$VeHjA*}7.owBI,\rY>l1BZsa>IH,>Hau},[2
    E>a@^_D-e{\JU;+AvJU7>'aT,+e{_~AE':WR##;OJxsMZO!o[We1$>eQz^oi$_R1$eOkO==<8^;p
    urXA2lsZ*1Bvo'}_ZPuU_ZV5rX],$>HRK#L!Xu*1Oura=Yj^lT]V#I}\LP5U'G,pz},pwrD+jX:C
    ZoY'Bp!=Kr^Fajse'w+3:ju$'S&y4~wIH'pZ'v{\rnGOsk]+-SL-pGnIdRC'~ji5_=;^i+o2!}@-
    #RrjvrY?5U<e~Y;oDi>j=Yi,!Xap7$e]m}G;nXsB}eGXG-e7Gp'*;7CZ1^AA\epe\Y)zJppXHD*^
    \rnc!=IH~_?V7+V{XOx*Bpl>N.)v1aRGn_5n}iOGv_?<zT?}_JJ$mRj3R1e$eO=5AvwM]HsU5H{x
    0BGIB:tr\1@^}ZA$rIB0!*Ba@YUE2\Z!hB;WzBGQ<E_]Z,1GX}lsp-z}'Yu$'wj-Q*K-Hk-]'}i+
    !x\H?2\2G*@JrluYBY#7x~Y5D:*Z<_,#$an-TY1;}<UDl$YH@Y>XIIi'JlQB]@'kQn3reeXRVap>
    {Q3VnsP:p#+u.xpCK;j#[B[BVR{XvXnD@\kZ'BmRp1.Ks}pG*@'}kR?@vBJP7_Uel'^5I<<GirVH
    OjpRj5EHl]k;Z}zQzJOpaV@~~Aa-x]TpCx>@XAXw%}pYECD]VjOpJR?R\e?;ZEa=X}$>e$Iv^H*_
    ei*v^x_3w$3E{*U]^zYWAx\-u31[v%5BJ2j~]Oj*}>!+A[pzT}2+vHBpeKIoUriBkT]2x-HC]?C,
    i1b@w\>v>\X,CHB>r}p?'5YxQnnnvE_^]ZBl=XpQRrm-pxEQwzpkH_R)w]E^BB'v(<Go\}>2n>nG
    >lwGZve@+^{Ar@n>3[DzOks]s'RIn*JC!['<Gse72{X'C~^&a'p!Z,s@K>OOvmv{jT$5s1[RIOzZ
    )Ax^>#Vl^&^{]*DZ!^prj_v2<1m-bOr]xLY3wrQ'xuzOrQa5jJ(pMD!suC[e@4UnA>y$awV7poKR
    DWl**}$E5Unvp>_[*n5zu_2E_Z5{zx>TX2Do?oUWRxR^a}53Dw?ovJBn-3~Hv_3I~j2U<OJ1>vvI
    GDz!eOBusir^^BV35^uow[IY{Eo-AzAevxj6/=G5n_5;CR;+[l+eD9Cl;2MMDK;7_\IKRe?RG;lT
    ,5wTZQ[*lx?Bz<*u~BZK$QKH9-GYn9noKJ0Kz\-xDw>-_?W'U;]BAD?Q=GWJ<1~Dpj+'1i2:dvQZ
    5Rx,ns!ZnI\-e(U5+GB\-_JI2BR,<V;-oO>oa2*wv-^DljRW1TY>jeWnelp]7mAl{mp'Rm^*<U!a
    oJcEY_vQD@Q}i]E+>]vB[O*-1u=_oUwJGDT4os!;2QYa-I1uRn$~z*InR^w]7v~z;pj>Xt\w7D_W
    x~0jAV~{<2wR|B1GODw~]HaX}N^[,R=$;Krm2}13<\m[1>BmR!EIn?-^X^m]<sev{H<$rQCB5mR]
    l2C=O\$a-+lKmOzI@BuU2@A5z2[\$vZ7[KqC<RjC'rj3}]sDupo+D,{3w{E'Y,^$:CG--,mxI?]u
    TYm'X{e@v#l@jl@rUQnTz=o,B-j=x{BKmrZYU\=\lan^JTDG{*+{z_!~5^zwv#O+K,?}Az#l{7D^
    UL2^5-\27=[*@GaGi,*03X'}m\_3$u<T}@X-VH_Vw'nC\Lx~ul"(iB+uu+EX7<z'T{*>v7+WzWAW
    Q?Q]IW{;$IzA^VrV~5$ju7-Aep'<$\[kYw<YI7<J}II7m}Wx_aOC/2Evzm]+'j#+wq,3QWV'U=om
    Ka;Xz3V'5R7_zR*BCX'=B1a{w;Yu*Z\}nXko1?)?j*Jp^l;D#m>(8<T2UGT!aOeZ[$~GI$\ll^Tj
    33'D}D*UK$OXx^v~r]UooRxHV3Hol'#}pG7^2J1zGc1rjD7UxC;^3Q\*nEoljQ,-Bpd]^~lT=opp
    xj]i<B\TlQ-{n$?z?T_@1}GR]*T}@WI'2A$io>l*lX7l1G<+nrK#5U!}}?wnRC{pZ'pEAr{VZ{lV
    $}\!\a12o>GAsE$QwpDeQQ!-BT>-7\ZB}[>CO$;x{7I3zsu!pslVjE=+pH5\v3Q=^=u*-X-u>mQp
    #Y'A_XI^~$Q>7Zn~rC[k'ewuVR@UxPz3=<rn}~YC]xcR$BEe1[Y9qj]-p5=2DjarmQ1GJZ$lp7~l
    3Xan*LE{j~IR>xxCK[QCi[mUlBDHZG!IIUQKAnw==!B\@eE~}u(iB*O;T@5xG@}JCJv^Bo*mCx~l
    BxDB';<\wx*m''>eKj$lXu{I+Xu1u$mA^^^]oG#;1O\p!az|~'W\3l>;=Us*~YOZU7uD\,o{VRXC
    ^Qrr;5-WqAaTEe}u$]QoCrUnClC$}K_B++pi_+j=a-_'r7pVm*H^?2_\Re7zJL!\wu,Yi2KTEHUH
    KA=ERKEs>j~al7wn3[QJnUnz_+5lzkarxQ\UKZ^pk3Tao2s~UYIa~,|#V2;C$mnoBuzjn2Ezs~O>
    5w7kQ_ovAGvTvJAOx[*=BIHv#3<jvT3aQ3-u1GzVZWxl=Yn'L2nvoK'xZI*z;VXv,%4rnzE_7I@7
    $AXC3KAlkVvvjTr*,z{^CK**~nlrCxnC+$jx;}rn'xuYCBavU+#=}Cvha1wEP!*iQLvauDG#supC
    #<zXo+>G^=Ie>W^sGH~zJZEA@7GmQ'pEoA~z@O'AmzoBjO]r,^YsGIe1xV3'GZO]A\k}Wpr<RHMU
    }oGUwJTTVoA.'xV'jQa\{}U1$J]kB^ECA57JQ$^Xa^\~G[$3BZH>?Ej{^KQi=pYXq<GeWYV^I]J]
    j2jDJJDJIv1$EG2wA7\ZUGR#1mw[3DVe?l!-w\PIXHBlK[>WwTZs$cVI_-T<YZ(Q5k=#nTr-Ae>!
    A*o_~_3!EJxvk3=,zs^gs>l@ovj~R1n35~7*Cw5[C^<=kD'QeTKww=B@+-3DVaW@u<QIlY_jBCA=
    Wv';^1lz:2C{>EI7?*^m-YkA{#H*D$z]Ql;QGx''DdC57n1ZliEk+'f;e~,GO}'<CIkkn],RG{r6
    ne;[mpZHR;li^+p}K>G1MOzQw&]~Dm4@Q}Y{1=a{UDs;A<pTCBHl7G{QjJKsVnG=K]s-HYv~HsQx
    YCx+'_Afiwj>=:V3*noW_[-^JGe[R;-z}<Wl~37#}T<751,U7V-=?W8-Q\@w^xW@x>~jJ\i,;RDJ
    \\>J\i$Du$G[XB;Q3E^D=2lOB1EWez1>'YEE?~WvuEaB_]Xm'$RxiWo9V5o\1H!]FkURnBXGXMbe
    sI][!I>l5IIB$>??$rX*2W\OH$Z>srwi5GJnTQ,VB1m{jDR$G~_<1=>on@~><p=~R^v}{;Tm]CeH
    I'!p2_O<xCA[#>QY{D,x7rxo<C$Q[*$(}HIZ\v]K)>lOjD9*CeQ,5v}_<xessQ+~Dv?9t|A7V_<R
    x]UeXptfORVeZXx$}p<Y^[;;QTE@3EI=jo3eHR*{>O!~]<\oJrsE.\3;_G2D~~=!xX1*ZDkxJ#A5
    vWnI!_rGV$55<1r'3V[eH3rB,7~jiv@X+Mejve!*+\]X[G,Z]Y4%31r~-];*>[x,k7Vmj~vJm>RU
    ~UZ7nUoaC'yMW[Up3DXV1!z7e1W2I[vBn-Ua6n}TBIlKUeZ2@ZRal#exxrpXncfo^rrW\'2\YJKi
    ]l?O33nGWHZ$e<T!>1uZpkmDBn^;-z]uEC*3]CezI2Qo#u>W{s@>xoim[?w^AYpeB+uxrI!nAX]1
    'eTCuWvY~5-7:=$+!ljwmC'{7s[wlZ-^k#,XTW{rT:~CY+dC*X*_knpeAjZodGD1o&7~xGvBFQmz
    -Z}v3IJUQNpoYo|=eKGY'?m:Ee=^?'IA#Vo+kH<#3}QCG$+lIJzBropX>pn2@BVC5n=p?1D$5J=H
    ;.8s;B_k,,Cgr+l;~jwYVmXOYCV-R,\e(2s-p3nDECZ5igUpaUDV7'Dons$D\Ig;EQui5+=~X12a
    Bm2H=5]e>OJ{[#r#7BA*j[Q~e;'Q?x@*YY2]]r>A{2,)lC7[%^WC]E{jOqJxF/^2V'j$+YZCejbl
    _<^YpC5kDoA$IlQpk{uIuns_w3Tg+<KosXQ#ZBp]wwC,$D[1Z+p?us+n[W\uV3lZ>[$1"Q<<HByl
    RVQGr><~^Ci)M!aKI?IxGE?X1iX[e[+Xw#,XoNn_23+eAKlz!Xe}KBF#DX<;R!j>}n,EEj'[ZT'M
    -${IY'a7r;}\B#3z!AJC}]o37}r{#<s+2DkwEBm^$Xrjm1?VC}kzB2Q*aE]^*;CzgDIw$*z~r.zj
    5KR'WE'eB7Aw>>5@JJ@'iI*XGeMH<~j=7_}iRj>gxD<O+=jQ:lE\Z{Xn3[l$G5a5Qme\{_u\QvvW
    nr--'*C!,wv,Y,;C]K1$'=aVR>C$=,kUJ-UOCE'lAZ<X'3woQCACjDli^oQ=ZYj5'S?7U\GnKj/*
    kw?1nX*ul=Bi,\p!DXu3rD\@+W*7wKe#5;'sC!U2I1Z+-<~^QCnzmDWn1v,<,+!k_7Og*C7z!X3$
    j\~[nV'!IsnzQ=G]>I~]q|Ypi\iIkJw7TWu[;,C[j$|'II{5Tn2HQjr$Q+z*o}]-jI}L5)YjJT},
    !>NCme2\!WJk7v]]V#1NYlX>HeX2j,*1ExA>pK^?1,<v<5?,@wr_XDQ'[2^;#T>wp-x[jlY[E?ws
    >-m;.z75syr'ZJTzl{QeHpWB5E)vjT$3v}XCuuBXl{xxX_VC_C_u,-K8xwWoE,o!jZ*$l_I5K'j[
    /pKr]2VRDBTC7}o_w?B3Rr{~Q,r>{G33$xmos2\RUaHAV#[>^T*X\>7i\*[;v_/Xoz}7{ACUYJ~Y
    +uB*a>;=]V,9zw-'Jr~QwaA~A[2mKVKJ+5uxVG2?T,GX#r}<pGmmXEWzwUeR(V@K_KC_G$3zwjo]
    7ks\??B$~@+PXUU=t!5nzXTA}37B!ia[I?I'=oi[rz\X?EjEm=[+JJ[',kXU@,e}JQ921HJoJKs'
    {7-AA;vE^;vC>,IIEnKEw>vopGuIHBuGU!vR}5!Vv$lX[sZwTpEEijpa_xJ~_k>p3lC'pYKpl2@0
    EHYv>Hx\e>\?]G-DoWGJG5}#$WYZY/irY@^7HCmQn*={aTQ2KzEOX$wjiA=^;+HTCT]3{@aE5~Rw
    7^PQaj;nC?QXX7OBj1$(p\>[ARip121^R_lj+{AHV>px,r!U)^XH*D'I}$EaG'3pYSs_>e{7{<O7
    Q<QXQaE2!=1{IixcGXuvjLGX$2Bs_*-QKjjpwm#X*OfHH~A[1BZ,r3^sr-,RQn1WE~VrZr,@pUEQ
    kOi1{EJ49r^~$ea<nsp[YYe\s]sa+@Bu{Z-vz~O@IjWpBrxU3]DX>T1Qw#$pk5nYpKXr7rB]!_!s
    #^kAsv=+jErZeA{s=HBwuKYB+BHGrjW_]emCkU7*lZ\Eo;_?>2*CZ*Vk;a]GVz<Ck$7Q;rRYsJYr
    xjIzJzHxe-X]IQXx^X}-I$onusT$pCkW!~Eli+B@]CXRv,xwAJaD5U$xW[EpJfaoQsGBrWaX{]UY
    \xo![v*IkX[Be3)-Dp]L]uR$g1p@'vlpB<^-\!\^i'sRuk+a!\G>#-IBYYox<-r@1aa$Dj*opCgC
    z!wrv;BO;{kC=ss3,_pc3=G5I<@sr*VJMEuTBI!aTxQZvK]XQw]n;SjT7rp*5p(L4EE+wQvlianK
    ]x$Z?TDX-M,YZG$;eOw,eO_[Q7E+_KolXHRT1#Y<[kBLL]u;[15z$wv<m-XBuEaHkeGxODJ_wEY}
    iC7_lk7HuHV!Q?erRj1oJH}@VG{o}TRwVsXn]8n^2s6},_wD2pp^lOA3R$E>ITm~}iJYHBuXQoJB
    Tp~\+eCCW_?I[J^Vm}+r!Vo/uv@DG-EZGG^ru."slAn1Ru]~^\j2=?Qq}jz5%]Je'2\1Jk.=YHz$
    rDD1X7KIr_WE^wXue2,_@Y;c&Q,2];1},w5Z!\[X[Ae5WY=,?H^$loAl!H$OD1BODwIX*]C>5g<E
    k#^mQOEn72rT;\'1pV,]KesVAoL*ZaC'R{sEGo@{U!OHo-{;XBjx[vG'x]1V'Gz)kaa}\v};#njC
    <el;Gx@G+'z^";O!{__,z-}R=AYGG8*oJ1.*Rz~^,jU*-+TuHX\vSxxUDl'avW5<>Oro+({''Z1A
    <s#*ow$}Qzm+$leBn+#'*~5>>!CGQnisTV5AR~'i]X4V;HR>UvBK\gmlQv+UZzG1jAseX>XI,;Q4
    ^KEQ?D{n[Z1^DT=n{AUG$3+IQl}[vT\V_\,QMo?13!plX^KJT.b,z>]r*z+BZU=_$}BO+D??+5#@
    TE3o<{EI=*OmV;_{-*JG@t][*^'22JI@xi<zOj{B@GR^elYY]'iB[H-{+'#A]Xok=,vImQ~''*:}
    87WY+*T}j]V!
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#@7KU.$]r_]@X^?C233e?e{Oj{$C@w-^2[fL1FrdpG*TA'z5%G?Vxv_-$sEzO}?rr=W[T-Ue
    v8<eXazxC[EfkQ'Be-e]iXa[zx^QI}VCX$sD72[lNW'#Zz1->qYI7\]YmB~a3[[3J<|9A9Apqk_A
    l3E;*\%~YGVv>v<g?$J2r><A2YV166H-r\;jKup}krGv7~*l[Q=3I7u_u}^X}W=eQ^1}XsO,w*o1
    V<!$\m?{C\2*!D~1#OI?<v)7nG*v-7mE$?j{v+<=HC$mCB]!=@}7]O^,aR_f=-}ni5#a8^~7aQ^r
    ^v*V-BVu*usBW={xxeo7xHX3yIjOr!v_;x&?QDCKAXC3a>ziUu;AxCr#_w=o2CJW=*EGU[Te#U;[
    ]Z}[ZRoJ5!6Z=}1UliV,IJ$xw1#s,{z72Jz-$5sY__[g_jBi?s]7VxTCQxJaGW3QD^QTY;V~J'_C
    s7n}<5Ux]nu@7-XBUvIld"?,<j~}W@?vBG-Y_zt;=U{a=5WGlDJ*+rQeK;xAe<H[jw7UB7]<}+=C
    pUC_^>7JD+l#zGj3xu$Cw@V2TZU-BQJ+=B{4"EkUZu{]JQZTOYA[[IE=VeHJenVjT\)+aYZwRT@p
    i{rl=\,g7Oo][XT!_C#-K5vl>RDjzG[[ess@$5VJ=HvACXTGlGSkXr~^zjU[piCzXr=v[#B[2jXx
    ->2C]A]pV3!2osmOaKsRw,\wHVHRsE!e5W_p_-pRxV+'\pafEK]$U'Du}A*uVN=RiA%5'nwj<uk|
    MlJ72l~DuEHuCvrv'eO==$~numH'_;v=![D]?w'Uo@5VnB>G>DOx,Du7[opAAEA^YQCa~'BX@!=C
    +r@p}7U2KUo1Zov\Ia^KB-$=>0]!5T#{OTY@wJW^I{E[ax}F-7ACm-n!<[R7i+AJs_~D}RoxUj3a
    )]Ii#=r3#]z@2TC?''iapV$,xA-7>Ar,iYmB]RpG'|O-+C)513?k}Z<xI5x[}QiO3C;|]jQD:wo<
    };*=uN>zK<DKXK\;V$7XR;oAap*X_~JDz,j#Js1u>kH{.OReTv_~1{'jRWXa[O^#,IeAmJvv@QxV
    Uo'VKVG{v$\D[6cC/31]UH}#_iH{1"r*]@:^Bnz^>A!'sA;u<n1*73sp!a^d,wE~O+e,73_1\s**
    earm\7-}-v$-)![T}skO,Axvl^sY#QV<#H^Bv[X]KRHR{qEEijV<=Rw$*ow^@>xs\a;VO!*T5J=k
    >*Yk\~vHZ^HLUCos~r-G;XX#@e?eRT\U_~ADTC!2JoA^J[#$/p!Dx5IVi?Tr!ieK[Z&oHR>mXp+(
    ~}m-=UXk3CX~GK<{ZXYkxH@O5Guof>x#s?*3jfwCal,;jpE[J~DO@pO#[Q=x#W}TZr:s;!CLi*^]
    *i<7A-nk~YI<7u^>pGT$p,#;=+U\sTR2LgD>_-7\<-*;Ox<T=om{$#lO]ZeUYi![xu]5oX@7n{3^
    i7,)aw+Z,E;!@t[]\]jXm_eKJx[J@,KV<USlYToQHEpPKX2-}v@xlBjBHepEDy^VZR;jG\mQ^w;7
    w@!eZlDien=J.gUa,x]UuQ:7xKvkjGU!eU}]B2@AR\@qL+DY@Vj-pkQuvKU<QDHjOQU[sxsWAvaD
    <Av]^m*;-T_57zZ-{5^l=}ZC7o*BX+<vALJ'=x[CJuBj]kJVXZHjDAg^~m^Q<TQYkY,zUY$;A3u7
    B<K1*<pz=TBj$\3e>zWGxX[~e?}e]Cz]?}s{,<sG;Q-w1WG^7*U*R*K/nRWauYi3;I{QSXBkuR~C
    ]+1GYuOX+>_Ax-jAA,CY?QQ!5:WEEEDll}Lcp%IQTDRGGv?e\V2-VAZYvuYKCJsGkWu+-X/}s\V?
    $-?~w>3^KEz!I"!]}J>{C'Ul2rQUj-wO;TGvJV+'JsZxvXVZ7eL*;}~<*Xam1]C\G<>V=Ujp#,m}
    #pKKvpRx{UT\-3E6Dn;$Bojw/7_',}}]K>\$uZUH<%7__DZ'~]p5UB_kJuzxGvqwY7kW_]!\{<^y
    !OGY_\xW<7\Jjx1#{RAAQ_+CsC^[B7Ue+,1!U=~^Hpa{>V?#bFW1QVcUvAka>X*;Y2~V}_@2l~5}
    sv--,Rjx_GY;_k]$-a_R1$k*T'Z=Biz2TQ>Ip_~{,yQ3lOTGBGY!{2RRHkVkx'D{uX?V2G:>qxmp
    R<-$a$<{>6|=Q$2e<+Zi,C}5@]j]spz<w@!UrK3ip3>B1s\2$mBlJQiXr\Z}e~QWwn3N"Hsl#OxK
    k\T}UYj=a^#CrU7V]YTVaXA\GowVW!HVHu^lupA7J+-eDGiwooR^}+_w}f]2,'5D?-5TXj;*eGD?
    >CV2@<N1H[KyR]oIdf2'vTqXV]l^;$p%-B[!O-Y_v2IVsD~$GoB;9,^Dxo2<jQps7a<Oi^;e,m=\
    746a[Y3}=vIe?'OmsO_Q!mR~Vo?3TJCplOJ*u7WzCEI+sHk's+315WA_lZ~25_],>^^25Q2ZsQGn
    }?VHHsUk-mBwpx@]u>l\_+m=kI[}OKQXr$2TG@aIwG!~7n@#{=Wu{JEuBIs{a7DZok+Oj-B]}_JW
    nm]!G[3V7w+lQ~aOOGV3EWYZDHZK1roZ<H<$}C'sYr1he*AsB-XVJDA@Ous]oQ_']Hu+yknj+}~w
    V=D^p>5s~[KjJ^lAuDDG+x#'<x1?>oK2!X7i\1E[T#^==^A{\Li<xCF'wau=,=Te-o\!D7WoJ]2,
    3]ssHYxD-HW~IZA*EB'p\{55[nDZQYn'@=RG_@Rr\vU,u@Xx},x%p+'?,vRCVsaj?V!v$]]m<Ev{
    >T,K_Guf!<D^e~pW6\'B*WCZ}Go}Ho]E!7\xT*~KmkTs7K$ZZ#|~_1D{\CETOz'okH5@}]vOwjY@
    nHY{,*knlrTiGNnr#W}pW,-UCYEjQB0'm<l?]$@'!V}{rH@7m@nl3uJ\A+s!V+sCrn}x<*u?O2w\
    #'n6J'<ZGdp+--'ZXBBQ1~A[?T<'5p*T!O)5EA?o$Rwl[!lljIiTvEVVvmCgvm<xDr'H=/#V[CI]
    5wrX^n_QaGe2=]rs3u\^poeme<TH[5a=iH9'e5{?B5;6GA>a7lm,AUXA73YC~HKWl<Usi<IHr]YR
    ]3JD'[k;d}>Yn4;<z5l2O~Qk5oGiGQ\_zVno>@)jrva*g2=u_f2pxiaGVWCGspa-V2wTT,3}+3Bk
    a1qo=IDp13$'OvvRoLe,7\Z<\+-oYA?oz27CXu5mV;W+^~,p{n4RIa}0A>1G_a\{JIk*Z}m;+5l[
    {In3{wE>~e{Ugg$soYQ?DalU{?KlTzjkr2R[sji6-CW;wU,zB1^+tG>p{=@@;DErjZQ]T+a}HEO*
    v7_ijX';W7iD~5<5Q!<jevB7[A-[,mIGo='a?jmC16^Z2Jr!$HiaW*:d$'>}jAs^2[;n<T}@DJVA
    ha_\Kxa]^sCzi3e+R_7D_@G^,p>JEwHCaC{ZG=l,$nD'3vHTpoyRm'Z@UD]/$CX*7a-+jmXnsAl!
    B+WO5+ok$,OKp{s#_QXJ_~U~vzlZjOwj:ARBxr{DT5wQzVQ_++RJCyE_mC-pDE[<usTHX+>HOmR@
    oDT_GV8#$E2ODAoQj,w'=Z5ppa3;n5U}<CwGsv@>CY+=_WnTz@7X-ID]jQkV]BBJh_#XvK<K*XxB
    p;*D?i^7H*u<omjiG)_ZaJ+A$Y_njnGI'1eO2w_Tv|>,XE\31;=*~ohTw@[JQ2#,O{7g:]G7nla[
    *O5A>Jz]HYj7m3__Jw'In|z!vm[{pID!@zY^*}[3TY^7oRi\!z~QiA{[+I]Q1J<5;{va+C#ar[B~
    $sWx^$#w=w@C{-isiVJGuve[j{+rm*E+[_Pe71C{op'W[$]VC[GO*-]\*W#*V7~jK{_X^QW,IuC^
    BOJXr]^JI<Zo+_$q\1U}QJlA!Dn@iIjvu]TC^+OY}DR!,Q-?2Gx-A>v37<x,5Q<umw9|3^CY!7Cr
    7E_KGwHn^-2l*>VD,e+@7#<oW^2X{Q@e#'H1^?nrdp,px>j#WO7mn[1IeBD#sEQrxv{jz+CVkIsl
    GHznlPaTn*mXv,Ho_s\DkrO5_T<v5Z7j,Z>xOKr25ie]-<Ja2E+Q3pf]}Pd5?{w5K1rsJjJjuYY=
    lwWs\=JV}GX[X=+sueGQm{Q2za{kCAQ$lCKBbe;1+RiDB~$vu*X$Kp$-R1@Z#K,uU8-UJK>U2eD-
    W@vR^s;{p]Rn*x'\XkmpvW;{DnD+H>RZR'Y8"@\RYHxa5EkDk\\W;}2Akx+^'lZCw_uWu#{5uCK-
    s@UT{2X7Ii$rRpX,_r{IrjRl>OH>+4<tmAQk%ZE#ZiaTKR$*DfkswX3z\p=ZT}?tJER={Q5K/:U[
    -G=e=w#U!JA]?{#ef|I~BG\=l'IFXs*7f~{5Q~Aaao3{~EUHnICmaq<DzCX*rx>n>5+R[jIx#W7>
    A+sup\C?D,jIv~}Gr^A_H^,Q1Z-CWIIoVRQn{5=I{unB-VhxD}<]Y{Y'>,$Y]'rHQXj-vKX?O,]A
    7ZHzT$Ax[iGm=Bno"!hiC}BQ,+U{l+YZ57V5eZ53GB<Yb=oQiDu=+*jJ,TwpXlH53_YKu^C*pD*1
    uIHzV=d{xp{oo?;!xl_<hE3x]wBm\M
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#i+XR[DH!Di,#a-_pVnu$bT=is!o;uOD*[8k7T[:JD"m''*}o;w[X^ZO/'kaBp;V$3^A,sZ]
    3}xvk=)_rPlwJ#*+[[o_n=['CW!Ul$HUlIH-BA=O#QET}7]3vTmh)DV>^f!$u![?ED7#YEp\?[k_
    Oi4ElC\Yw=$=n2Enr2TAEz_|k,Ap8V4Bn!W@'+\vjm?_ZzWA]@sK+mp='_oVD+}$}[oR3,#^*1X^
    1s#t]jJTFN[ZOBuV_p9[{O='oBC4VLcAlz!@aR$jw*+lHH7O$nrKo}2-UZ<Ev1leK~#AVB+oR>Sp
    Qeu@U!B,z1\\wjItiw,zW]Gu,$+oJn@mSjo5wQQR3qZ=HrR$nGVrUv*W]*{X-O<Rn<.P{+_#5{m,
    iem-[l2'$}iBl@O,!5'5Y]knCHp\osTKhvHDvTY{ZO+z[Xe+-0EYYQ}BspT-pu-A<T$?[u*<pEIC
    @vU=Qa+Q$k$XX?7!OmKe-v0DkZJQa2T8B+*lxCUa._v<l!E{lCHomMkUvJ]\^_v~Q]$CID+5?C=u
    3op=Y>72vaiv!^?_3~#XBW?Q~lm}X[rEw{+pY^E1#pApUU14c=Y[2}^Q+:x3lj<SBi3*b$s*QVG$
    [Z5uCav{]kn{viRWx*jx[Y-I[H}+O-e_v)NO'jjp?\GYo@\Vep?{B?^EwHVzIR=DRjY<'+=(u'Q=
    X-Cr1<*TsI}Q?<pEl-<a}N}@R$=ZwJj1\o{e>A)z)!}$1![=;^OAD';mwH_@szRCBQro$52K]EAQ
    AswB<'euClk5poG_]5v#*NJGsXsrQ~vK_J7J>Z@7Zud5u~jqEs--=+Or[vr?*1WZ5p>Zu]>\WC1n
    0{>Tn@*@=+oooiG^iNl!J@2OUW~=Y3oQC@9D1DXuj'7$A'{7ekx5s#ICD]G0zJKDP};o~*'}?[2-
    5Y]Drm+H[)esuxl+;k|Wv{@o.R,JH,vp7ae7<^1]C&5i^D~,oJD#[7yHaG$2sr#{]Ez'UO[URO!J
    xAKjReR,,DVxemE]RiDlrjR5n~C;GUJ<vwu:]DD2?_BI~'UEQo#ook<;vI$JwOwKh?Ao~X$]<Z=w
    BkozBu5ZO=we{mzY?[z1>l~~~C>^=uI{T;'ZQK]OY"[T~KY'uCoLKEOrbRxG.JGoT7K3HlT1k'=+
    $2rO-QOp1$Vu^A^2BsK<oCu,rcK5KHG2C]VvWw',OlK5,1ZC\^Jt59KX\T'TI]Ao5O{lZ-'$<zU7
    !;+1GU%=_vp~7[U<U-*iX-B5e{xl-C{5,J!sBA1j=o_iU[~,G#7-1@kX,_l2BswsQ~v*z;@#Uu!D
    <u55iD<_#ZTA[Rz^3Qz7Emr6X,j=pvOa27a<VnTTs-H#GsT\Oo7oH,X7*<-IRB_K>AJ\DHOBwV]s
    ,;VH7{+;E>\ef2,e2o\TojX];],r;L'aV3fRamK,{E]^sInQZRQBJ;*jHv?1)x2WlxUQa1IOo's5
    Z#<R-Xp3x}>v=g5Jura<[p,-In;5-DfQ{u;Gajr5E+apx7~^3]$l{JzAv2UE-UmoAwe3>XHRooKI
    Y=W'r\,x3jHekOT=\?K5E'BOOr}XE#]'!jE6H{_*GT;[JT$rvGuT,HuVvKJ=(1sX;jw*T_<lv}{'
    an]7W:ivG^RhYjuu?*!}^moJ~GZ#pO>_!oW=Dw^rV2[]wOBT[g\uJsv~5z>pV\w+OCk>VTs;rpb^
    AJ*cD!-upaj#4Bz\O!=+odQi{*#X1\}Hr*w-KDeiOK$$,pr}!+cI<j}_@VphBw'KJQ'3_X^'x2@B
    =-_V>*H1F@,ZJG~TT2G~ExnaQlUD?*HKWm7T1ZeHo;n!='iro{UWTZL35v}fB8~Tn3GKH@xlE[Hp
    G+^~3V,rg1QYwwDOQ{rqO+-re]aB'[!_O.(k,TkQ3>$27sDD]~\vwnZ2G'm7wUD?'<+3BX1W<xzU
    BCm$'Rs(OK5=JUI{jXORk-x<7!DWjw7R"eOA!nT5GGTe[\Ee1z2nRkB<x^vOTX*5J+Q5I3^mT_Vi
    -WOivS+>vX\n@;wr-v9,eDR[G]?Wwv,i7Uk;sOU>Eir@GrG<H}rk$7vGU*ZC@veeE-jE'IJ'D=Q1
    +XCC#I7x{3}B*;Btoaji]B=TkO'H!Q=v,7I<RHJ\0GE?z3ev[J$xWJ[W]HXw#15[UWrpR5i]eDWe
    5BCA#w=aK~<_o$E~Ev_^aYrAOip2[wzz,~X{~jO<?clV^lU}"a-{GuR{[uw4yUY}o#$vll+Cj{}"
    xwZnB+z;
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#Ep@W5*A_lw2ZPY>x$$X5l1QUVaXZrjB#[.Q>$[I;{Vh<5K?@QT=75Kj7si!JTH$aUC76=lG
    G*_;+<'k$_rPlwJ#*+[[o_n=['CW!Ul$HUlIH-BA=O#QET}7]3vTmhmHnj1{<*<<YuW}R^CeW3CP
    Uwe[V,OlN3,$7Sit{w}x2l,uW[mkH>Wx,j3!Z_HW}+KK)-7Kp=QX^V3KlwC?D[.QzARa<*{:<lTK
    RomkU,~#]Ri1-eQ_pZzVin2}mX;Rb#$ZR'?=^)y7aG;I]jv'5x[*o=mx+'\~VlWtiA2592,BIQ^_
    BQGp;p#XaxZe*#YGuzDW!\=~n,xirp+O-=@WGZ>Owx^7?Q#**]@$v{Xjipspk!=}O;x$'#R327p3
    m|&\"r;U=h9e{R]Uz}Z,^?@v]5=j@DZ4\X5p'jIYt&?pXTNo^n;cR>lO$W]R-xjVajT?UvWDr,C^
    B5zxP{_][;GBw*#Yps$o$.lml#[YZ>Gk*QPjC{xp>x5}r?;Zl*]C=_p#5Q-Vn@=u]Vo<AA<HQ>2M
    "o?K-HT{Q3>_oQX-z+R?vuQ?QVfWv3!Z\rT[@$TxIukDtIUWD{+oYs{*Xjn~!GVBlE>\r@R@CsDi
    -3wU<oTD=*Av{k7rs^*piLAAjn1-{#rlK!Wp*[7TElyw-n~BrR{KnE=RBVosm=pR_#wRD?QJ_jYi
    $j}aUo*DQD>VCz[6OxHA[A[2#w=nFzQBrUY#!>[n\[E-A'C]{?a~ILIJ\sT,kDD3x]OOVY+R;B,v
    ,^X[iVB\KDe]iV9#zp_G5[;]iXojQHY}l!rE'ip"s2Yi\V_E7A*@55=TB~B7!w{K-5k_rs<kK\u>
    7mH{Ir~TEna'YvV7:!'{3\We\,[+j0xpx3->*3ZR2jD+K^E(R~7#V}Vm<HZnW}vRKUhe;Z+4STUj
    <\naV=i-Qi{{Os~x@}vX1nxp$E$$!XjlJeWZR$3V5QE\'xiRCsBQ>>}Densx$WwVorQj_+RG>@]i
    Z#-X,rm!>&xE@je}K;Y+Jl!-Ru~7[{*uH>JHG5qB{wZ4'uKR}5#pA=TQE*XT-67ax^Hrw};1E\1H
    }Z}GA?'RRi+a'2KXz'u[>]oWA;@UI*Y52x~5D3$J,zW]OxC[Z'gDT<?r#u\q4]-7ek1\lF'3mXH[
    \V_Y+j\K,-lBx*BwU$='arTBwoKE1$H_l_?DwHFdC#K*vJnI'0YupmE!]rs+jCc0.DBYi5a<,HY+
    5y]CUZAI\sZB?kA}=V8hW7?>ea=lE7pm~Ts]:]T!K<ldl$]7<>Z>I@Xu$$xOm>rjr=3Y|TB5-Y[>
    e2_pYjp*l~Bp]w1wYI;<}Z5+xz=_V=rsoa_Iz>YJCG{Wk1eR!7;lU{s$CVsmwvJ$W}kUk9[I<7H_
    Ren1Aj_eRC*?HmE*WXeHBoaT]>LIJ{mD-Kep<j\cTQ{;'pzl;$Az|_oTuj*LOrv{<BxG_~en?p!m
    Z1O]&H<JQl@x1^WX^?C>-sxKl,2UHC-\!pZI]sYDo^j@m43<_W6C5?#Gv!W_>XZVC3Da}'_uABu?
    B#'~]*]|j3,C@nIw:z>KKO;lB,oV=Y}'i)Enr{hH=,^TRu;Hw*[=?GET]XQ:]J\X*3}uEYk+,#Am
    nj-B)'XZ;'B,7alGIBao[#Rir#]!#$<[V[~{BrvDk\O<,I7_e=X~DOKTv62Y[By$OJrnvRAzma[-
    OeE1DUr5xVJ]x>T'J^{~l=uetoCkV-*U'xZJA;r^['[XeDQ~J<Bz^p]2+mG2Ou'oTjz=iO'[][BC
    s7UuwP55-k-x]{@7o[a^\v_]UmmQ[!1{DYAq[7}=,H!5>l_po;ZT2{s,*_5{C+I$%r@rzj5\izr_
    <<+{2l=meQ\'2H<DnG3v,:}w;u\Un[_~<7u1ux7pmQwX*,'CVv)'z5?G<[=r73Iyt?e5,3to@uJ=
    Za\-p{7ti,2;ZD;m!5iCW^Evl3G$B2Uj?O{Gb/\K!>$6_;ZRBWpe}expQ3u5dHxzKeu$U7{E\2na
    {;e~uYoxY{o=EGsE<<$CV!C-=Oao-[n*^_D~Ku}[COxeYpe$U'@H$uVkR\#XHvdur=1Dev=jER@?
    >3Um_W*UA=ZBOwJ17?Jzea2He^'Oa*X?$7?r6~$1z!aZ?DA=}]zA~V>VIoo~x>DvArwe?5_><+\W
    3V7l[;CEz,\S3p!^E7A!@z^7\-jpABWK*z$I'l$I2$TJIk-xMCs}T%D\Z'XsV>~RQJREj>,saTU<
    -[v*<!p@Xkanv~6cU=AY\}X5Aew_i<VY<s@wWUoiWln5Fk[#\2]?r5H1v^F$$_VV-_5GuYsPT<-x
    [5mA_]J*K_jORZ5wBZ27E>[lu],G{]H1}jQk;-Ts,$IZk'oI~+BiE*11aCKp~G$R5>!E;TnUW^<^
    5x!$z+$A1InTAQX!H,w[j+K}w]wCxl>>,or!SOYr}Y>1-na~x4v~7E7saZ/rEZV-5U'^Tev+UE_5
    m{up_UCZGm-OERVar[2z>\_7R\m~*GV*2XH=Hv@[pl5pL1x3WuxoKr<]!ei-r=Ju#YTGvvD{15X<
    !j+Io<nw!=H^!DiA?a'J?xe1M{aRU^JGWQ9p@aw2rC#[1;rR>65KTmYEI<E[
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#fu\GKwsVw>,pIF\o#_-'O~fj3m{JD?E[)3Y)Di\?(H['Z#V_T$hTB-}RU_O"?o}['~Uvo*n
    ]-nXuz3C[EfkQ'Be-e]iXa[zx^QI}VCX$sD72[lNW'#Zz1->qYI7ppYmB~a3[[3J<|9A9ApA]K_-
    <?s\;UoGwaoJevH2koDQVB9Z]+XZE<YsuXTxmI!i\XC=3I_93psA*}He7;*eXBY^x57u.s2'#rQA
    W~+OBsh#YRp{ta5U<+IW![T@x+x{,~DZ^WVip~wDTBTUHknEEz{J~HTA#5D@+G<akXe*i#>B_ba{
    17=*A_=CHYoZvE$e=oB;2w-\7r"ajjkBI!+N+lr-~T{_'{siRKYozrB~|wXjY}?ZYSmji\lI{{\{
    e~U<sQ@Uwe{ezx.xx+?'}Vvwek''zH~Qk]s$*[@=iO-|k9B=~z!\RY}lH\T}pYHsR*r=oBwQiBH$
    1pE/=AER>n;#!Q;w\?_<lpH@i*wDG}HBz12-,O1UipCKwoaX]71oXE=j~_[5wj!vWV2j{w_'YTH2
    o,WACi+u_CT#2owDG*ZIaGe3E(KTr=^i31REZX/ZD=d"C-!$^dC]\k>Dt#>Q7:#TQT#Vf4]]5T#1
    X-'+AeIiQx$l?HxaD-oJV7tRo2T93G2}xrCw$s[eE$;WX,v2;z>#*cE;z2rYeW'=73pU+CH[n+u-
    JKyl~$mW\[wmBpGY;2@aYVY*R>W'OCs>Ez\GIn<%#X+oBlOo_V<{]MCZAET__ZAj[T+[oT^>UuOU
    o=LUn!}(C}?XB<=}zJ$R>UT3hn^Zl=>pEVI];zDD{A,uRgIJ*#}z-~XzvnViVA<Q*Z1>n<6mH<2A
    s#CFojDGD;{oIx[O1[\Vnn*QJ>Cux51RB_eOa[^[o5>!-C^\WxCGB][7-<v[]eTWB\@32Tw-6AxU
    K};Uv$Uz_zxm2n_zp[DHrEqp\{{\2CI'65Jo^nBET7{^HC9A=IW}U$lO$#x,\G^(jaE-Bvs!NeXT
    \DjuZUAEDOK_\+^x=klr5ouY>YxImH+$Z^;xA;EuRQ?]JoQB2==sljHv$~XK[15x{ovaBaRrXG]s
    x5#d,n,m{HmahO3Z^7ux<~AlRY-DGG{=T{s$oO!BDwp2<*IWKVx3;2z?'d]x=}j}1AYiO#B-pw&[
    }}lCC=j!HnxvFIJuo2BEGCz-!!s]@=^+nE8l6^kZk5j{!5pz[=~R*uY2CE2Waus|r@7$wGm;J<
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#TwvVbv>3G^1WX,$@5E<HwWAw~G>TjKA9b}e/$@_Y9<}R+@+XTjUuoc1uDlmxY$_he?7[wD@
    sqC|z3C[EfkQ'Be-e]iXa[zx^QI}VCX$sD72[lNW'#Zz1->qYIljvY\oyjJD!l>p}aDV~F6IZVou
    XW]6aHK'}m1mC*R}VuC[?C>Ca<}31-$2lKYrCsIIa>C@>{;A]w@u?R[?]\1\h!=+-JLEU'V7)v4Y
    ARKiT^iEv+?0<Hek>-a~7WzRB5l{a[D<!_(HAW3KwnJUazW]!H+Ekr{7'W7zd$B1WWoZe*37DZlp
    <D}ikX'_C=!~oN+s?,[2D]7usQJ+KTavW{\;!U21IU3>x=1,+$25u1^H;OC5-,!^_}z7i17uB2]3
    z=@'R](2pBu\IAsmjwDO?wj$+}73Qs{fnv2rKT,K{o<Y>EKzYuK[<GYxs}$2D${]a,rXXl7ru<Qu
    l~a=JDppj>rY{lGG}l~QPI=@Qc%m^-H}J1E-L5T1m$YYAEUrZUC<?0,~EV>_Ia<[O~=JvnEzjA#{
    W^v5Yur,Xw|Ja{Rn(_7#TP<>1#~{RR#nRV/[Y5,-Iea\1,ex\rZ$K2Gvk=ikjZ{wlm~K[a36K\Y*
    r'7v:Q'TDi,;Ospx5RQ!m}=?'zWRi$2jZ;7XG55olP;x$'r#[\E![l7Gl2aY\aQ[i@kAp-R<GHRC
    {u$*>l_DjB.^,|-sEzWjk2ZaKo4!BXpa<-!2=Xo!7Qk]{\elkJ]g=_?Z-T>Z,D>\m^RoCzJn[*+=
    pk>KYGnvNZ'uvk]|]^5vIR@Jp]2j<7s~%:[;+sCDTGu}X5uAX1'TX@r}GnUp]H-=,IoImmuU$ziv
    an-[?>rv<$,[OEaQ@pMYw^\*KuGEev?&LD*rAZ<^2mTO?R2^$~G-auBACYaTO3juH1XVX^wz28i]
    $s@w@1TR!zKC{O@ex$ln-DC{jeH,>n-Ips5rJOkX;Olw{31uop[\*DVk*@ihHE\-p@2=TRjA}JZ#
    _>D>GZ5ID9v^uoel\m{ElwD;7XrJYGY-r!#ARlyBD*E;Y#'RIv\<Cj>E]p+-znow<TClK!X.5T;;
    X>lr^*TelAu;N}]>YkU7pBs[~AsXkb=DQ_N?Y$kW*^AgMGlk#Rk\Xq=*]B-,{BGBRDjKuur,<-&o
    Z>kavaDmA}OGp@^9D=T]_*CRI}a1FBIE_E<^HG5<]zB]z)Tpa}I!wGB6p~YVgzToEz{7$WA3#<rE
    CzMwDBV9RCQ;wI~}i=VTg9j+s!n-1kjuZ\3{3kYmY[C\GAuH!7(+Erv%7ErYjZmo-5En}rW=1rZp
    ?v;55az$k<JEy$;5Yyt&}V2{<}K[pXZ7Ck$QOeCjf-AYv35ZX7~5>e^$3,RZ'CR2D/>-1{!-\]rA
    pk*Wmnr_2sHH'<ZTz2@<BmG1SK+'5za[of|~TmH:Xzj~dv]1Oz.D{B#^>p?ERVZGEzTGUxBEXI2F
    o!T_=WU,p\!W{=<[D*I;BnR~(B3oO#Bs2Bx7{t\~vGxjVeoIQ*Xr@Q5TE7MD+A,+-_pYE7~+R_w#
    ,KxIaXX/9;{=WpK~og1JUW91~QX7k\AeQp5{xrX}!Az_@xpzE\nwO!GviD]=?=+aalXxv\[bde3p
    Z-sQiD!>-rI$,.CuDpz#l[eZm{(CkaYue}K\~E#!r?#'?n!>{x53[U~]>EumBA#y\}H<^pnw=#5O
    ;5XRzO3],~XrBX=>0e~Y2P^W*J}vo=S;Tu7Q@uA@rn7oinrk*WQR#R7eiUp'B?,#DC~o:iE_w**3
    C{O}zKU!O{{{,Y($2UT~1$R\$-2eVDVBkWnuX_2e]pj@-D<<[;n?Hun$>aJ;=}lR#WYj*ZZ{^In>
    $m>s3YV=WXeTA>pAwpxx3EQqSp7^rR!Qv']IKOuD?YYBo[_+j}$QH{'5*nw{sl@1!7}_vm-ZX\xO
    @1wVO7_z,7R\j<$p-YWoUsVX=laBDK=$Kl$D>lW71em^*Rjp}zGk7m]>Cz{A;z=Q?7$Z2u}~B]]2
    \?UK1[GWZU[?*;Oi}~l3HkoJo#RVn|'{QmlwB5zpJsj,uE++'xA5XUYHGzUY],s#rk8jADGwOH3R
    ={*+\X!El<U?[IBwaT~^rIG#v7HUOvR&Epw_JaJzO][[5X<Gz2V,Q]GAxDn#>w1j2s_mm^mEG?BV
    -_lk$ZaTDY^+]Hv]~jk+v_jTOa,KbQ1m]Y%y,3{vfMACO_I>=W\A!$g%%>rOv'iGxPK9GkV?onV1
    I>K\41]JW'+Ka&<^WXi1W^sK'kjQE!rn\O}WJ#$9xn~*R2rm*<+E!=pn~G=lEzx#G+O2%%dd7eGz
    'Ov\,5uKsjp{-aH\z'_kG?e{r^$<Wr*++G^'{'?Jx{CDy#a3]|!TJeG^kQUlB-4Zja[71zpE_?]a
    7okGrZ]5R*2CIpHb6Vuo>p;;AIXUxIZnKRX<XEeo$C5nX?*>l<e;a/{zOR^#JzpK\pCQlYsnXw]:
    [pR]1Dr3V'U?}@a-p}+pCAxZ[I[IUDinCT{~@n=u-B[=kXQZWpk'*Qz[}<YmBAu}xE\WdxQaw7uC
    @E7,unDkHV,#-=3!D@nQi_KpRav-pjM1=Y5R~H,W\]ru1nJH1,*3n@Y_5lTCiVu3s\Ilv3J=KuAR
    eJ>k-e5Y[r7J5Dwa^]a*#72T=?Ix[Y-zm,TEO3{U7;?>_^_u15H^3m2-RYnbEK1<Er*KK]$rC#O\
    )i<2nlD\Bu]2\mY+@6<*Yo/mU+Gq|BO>VVR'217FnnEm^OQR}nWmcDI2I]]~D]Us@zGo#mz'H^3n
    ~xkTl-vYImwK#GD+_tC=!^v>U-5\5i(/wznwU=kj|Vz$_j5?^8C'-Y3A~GnEQvEe\w_pA{wD57pB
    u@GB<]Rz\aImTe}~DX*vTZ#5w>$AX?;pQ3v,^mjn;EI5s},A-HJ\Rp7I1xQ$BQ)f!Gl=rAD[=3vJ
    C[jK;8r!<w0[>5n7v1u^=a2B;!l3U7K-5aRY_~v-Lr]AG'{H@<Azz;HDa;1$D'Y,kGi7koskIs!e
    ui}o''![o'2^IX<av{EGE-o~Rp<BrQ5$Y{--_n5wW&x{Z,X>{vfvHT?zXx,,rp[ElT@R'{[R5Q#,
    'KYVQ[\!97wRu]CIRe+3IwCKGQ?$zvuCl0NsHW5qe}iu(2xA}QaAZs2@KJ<1TJneaR>~oU-Aw<Ij
    r<+xnjiKzYJ=3ipO@k\7x.s$HXsE1ppA3TQC-H]~5^TY!Y'kw?:HsB2ZCkDxEZW\2d2D_TIeT@u_
    ~B7#1{^-KXzme~v2{Ak(R?EWZ]2U,Lkaw#_C;5@-{;7+@GpiVwg5_CZ0B{H^iA1@s*m~DlZz_=[e
    n_,DX]QioC[+'KXIRvYZeulo{_JvQXGHjCks&]!$@5];A^XQ1>p,G?=alTe@VBQoJ[<!E?>2E{nA
    wu7^mAUEosoGx/i<UB*HI?JD\rW+-peQr,kX+]dIw]r]^Hj:?wj'j=EvGKKm#=mHzrn=_1p^C@'o
    ;QvTQA~O,}_3n-3,I#U@UznvY+a-IxsElT}2^omXTT5^j3z2GVO1(o5Z2SZeXpOanJexl[K<'#s@
    Jx\m;@S=jr1p$s\@w-e#DE;lZvx2Vlo[U<>BUXZzQH?UG!?Cs;>EevY?=XZ\m+pR<^*V+un}A_5Y
    e]afI=lCoaHwInWULzjXn3eww>XYTIzj'z{ue1[XZ!UuI~l[1CuQ?1.vkKWsQ2QA]z*\#$VA<JO@
    1>z4vavJvW-CYlQvx+JA][\J$,+^UjsuIZ^D$o@~>{v7?IDT+UZ2XD,*))o'mZ.iQxK@\AJnpE@G
    sj''x5W2D\+EKv]V+W\SEW[$#BGnz'$iGR>]'sIZ,~~7TYD_42^>XVuEs\e,o,C~mEaV'*Ia@_^E
    pn^!Gk]DWsBBGJ5]D*R,k#a=a'J]]p#'reW!]&J'}[_]IoeBu\vwHXL[e@V7n]\>r$!z,Z[Z1^E1
    znY]TrejXJDX=UZ&;VU$zA]k$<D\T>AQQO!O3a{er{!UJ+==Ev<>K>xOe|pGZ{v_k',W@H+XH}O?
    oIHTVmwBJ^,<G#,+InU{zDCDVB=e#\Q5-]QV>*6?*K~YppA}-~pC;}_Qn3n#}[>$UDngslW'#l@~
    };^r{vG'*kAv=v'_}<v[{5s_}AZV+lB_*[==Pe*o\R}e#WU{!e>Cs_~_K=]s@7E^J3YHATx=\~+}
    ^[?>CsETwp91TeHQ<=]1aGRJrJCf{_kO+-Oj}AKCI!HT%RzoU}eu^osH\To_TuT^5^iR>Xoeuh~*
    Q3Ho1A_RB^-','6E$vWBKQBeZwj!{]JzP;Eaz*vVs[Zzso~;#5*zT\_Isgzal5U[C'5*m]m5nRW{
    {$o>ZRMCI7*1Di;9}m;k;*-2TBVBCuA}pp,uax[]Tl}+IZIlK$J$FE{7nGEK=eZR1+OuQ25V'1KO
    G_]X]Sru7$~*@[>HZDkaVs_]k;1@C^x2;JTXUxOZ1zvI1@Z-ZV#QZJjWTJ^@+>*'IozBYUW+s+{,
    #,HI@}AnBDVsIuE#j^EksT0#To3YumEL)=K]Xu*D;U,;+naHu=\*~K'a2c_3pmgxrO7KOw]TTR_k
    Y1V=n@2n\]jp7!_mBGI?xE#s}5x@O;x$'_X-,}xHGkT]eBDviHDVtl+UHJDEB*~H$\slWlE5Vcvv
    Q~PGRn7r+KKE_InVZ[#_O1-z]],~=2_E]We;,U=1l$HY?<+WU7]HErlOxW$kC32c;Y[1TUe@;'vW
    \Gz$DRm2Wo;<Hx-Aw1;wYV%8PR~Hv,j]wzn}lTo;V!'=l+z\[}+-GWHDIKClTQ*]B[{*ls\rCQCK
    H7~$@!'VU3Rjw^jG,Ee3-Br{eC;Hm&:X,$]^$@U#RRE#+-lT\[7_Jz\]YEQw^}CxA<$-BD3>TIli
    A!zvwrXHI[3Ea]ig1<WwtJ{[=[]w~[\*3x?uXBQE{*Y#GC,#pD*^'#lqN{I#I0=A5uA=CTr-l,^]
    j\pl+[vQz}j^l'1}vr{G7snTVVns\YjD@X;\$KpzjDQR<H11njT{lHjA\Y3HW\4n{Hz,$\W%EOQ-
    7OU[;R]jua\GDUm~<[<GvC<3)T,T+9jAB-GT@@@enBUaw3UDeZ5#X,>lT<pW}_jo<RYDDsJs;e@+
    1]B^1EuOimpU>m=-CV^]rlZ7O$2IpaBWXsoRIO2o~D^{]rz?!p;rIG7a{:[;ep$#e;1,a}:Op?}i
    [!WV$JDo,;CB}rm,XOB[?+J7ee=R>z1[v+pbCo0tue^^KTBxl7@aX_eHzv-n5-T,ZjwY?Vp$v}ZY
    FDI~=wX^kRJ^pRt!Tmp*JA>kGka3-wox$_?}Q<\N7kY;AY}1UE=
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#vv$B^viT-_1QXDj]vTapg]iOQk<pBVZ[[I;l>="7*JR,xC'g2VBuT[#TF$@~;c?T2['m5*X
    YCJq$--s~{BBY6+1$'Q,AmOoXA31,['>Kj^-1V-]3]_7[{j'?zs?vm~-~JVhI_\1E$;uvvG[,uj\
    [5=oHonU=WF|d[ZBBg''w7Z17;x,u>]koO\|wUer]]Qk@=#oE~CoQX[_}Xe*y}ysm<p[*oChCwA5
    e;uvw.OO\?*<Cm?X@7HnO2TUo-i5orzjax9)=zz^}^pwEvV'X$V$}#{Dzr>HzT+[@<JCvhnD~<nj
    k~a=uGErW1Gmae3Ro'HwrX0(^rxzl_'>na+OCOH@!>XZ>D>ZA1u\IiK]~{{}!E;luUJ3G-Z5?,xI
    JOApUTo=je5TOa'J]~D'=W^H)plWB6}]3D)1{j\Vn;@iA*W}22@>1l-=l-H#>\v}r5<\}{a*5mDk
    B];Yn}}GVm@@51K,Z]DN$u<_eOOrXsm5q]3{H,o{QQ~CA2elJGl~G?RQQn[35V,Civ$n1uYjZIzC
    [!$[GYo+>1E_}xJ<JBH;}Ywz=*nsz\zkD?*BUDap=}T'*p]B<^aQO(]O}?~*#B$|RC<u^sUnGIev
    \~~=o;z-D!1?Y!Rn%;Ra}"gYJxW}$Bep#HE|31OAI>=r{BKrGCG,7*Xui'VVrGesQje*se1Z;ls[
    5>^=ZrU@zK+oUB']5TA<O?~577R#|aeTXaR#!Q}zoU12s8<-\\1;J?Q7Q=rBWUBVxA+AQA}}V{<T
    EKj:Y>K>@xe'_X$]?GsYn'Jk!'K@@w6faR1[?\a'rn]si7a5s{[[['+\q>ovi[!X3@C_!>{I&usU
    _r2xsRVruCI1-R\vVji,QI@pA41Q*H2v*[@_a1'rCxsCQw5a-UzK@@EJOJaOmn7u>nV{z>,[+[;=
    AQDQpUlRi#Ar=Je$u?B$=JGasuUGUJr[spvaJ@QY3](Q_dJj=^lJOK\51vv\Viz[}Tu}DnpeiIEm
    ~ztV~+kZ-eDDo[Aog2vu<:GIO+C}lDhx}o{t,vvWxU_l\WZ-'[?Eh^I\jG{Goj)$L+]'\lBA#T=J
    m%"\vYm=EoD^u;}j}AoZlK{Ia_+<VvjyU]{kn[>T,~+]Y!5IqiTVUt^TJ\p>[^$3<Wx{U77*IY1E
    $?Ysi~t8hm,W$YGi@~7nmqH1~^#+7lYij$e;K?s{_s<>,$*;GwN,=YAvXp}1^wV'w,=7JUWkV13U
    n_jDK[BD'OUaE\v*P1CO5*+V^OI~j+H[B=@Q,@x\5_@~r^KJ[}beCA'H57!'v1X]e~!ueHEuz3OL
    +U*X]j2DgzB?Ak[<VrH^YjIIOYOWKrOK<p5=n|QeKaUlsej,Z3P|:j!nG=*De2}z{[iG^Qv{#lex
    s<7m1uOoij1Q<Sz]{5C+O@'KC@eW^2wr!Wm'AoUxe?I-,K-N^KU\xpjk7-~7,n{A3BQiE&$^E~Tr
    *}@XmCQIHv\xi2A}-HY5r\-E#x]2z^pQk<%;\ReNw\EogsV$DJ$[pH7a]\DE#52z'Qi2O'/nj{}g
    $#sC^wYADw+a{AVim_U=mr[Es\-=S[$ArUjvHAeO#\nJJom7<VQz7rDrz+{oVR?A\PRx{^HoAu\R
    nRH'wZvWAAX=euVlCmKoDQC=]ww>n7^GwCN{wlZ-1,CWz~Ow7sJ!o~5iEn1#oa^[G<@*+ZW.pT;\
    >DmAA=#rB?E$pH<R6:)wUrH5jJ3YDa?T,vV&AwE@\1_3rwI]rj=YNo2\lfw'-?3o$[A51_Zl{{A_
    ;Z>OewjHGk+5{oB@mYl+CV*^I1o<@KHo5rxi>}m$^vlsI^5AVu1{@2<I]*!O1Q?HSjRQ]tOB#TO(
    f_q_iUuj?Z=RiUUQmr?-DX;laaZ.fI\iO#Up~EuDJQGG+H9#zB]B\<^1[T}7&eY@Q,ekr,d5I3je
    +el$;@kR}w^f0BiTXY+1-A^lp^<s!1BoHr3Ku6u=[}O*?\[>CjsO,Qz^z^K'T]7w[nT*z}du=D<W
    U-Q*#E['1x7IX!z;lJWwpA#w<DOk[V$!x*o*wQ~$aE#'^'B@oW$YRTU=xou=[7-*yZU$;pr!x]1T
    7zHlzYeR;jz>zXnRp+D]<Nr[HeFF_?-a^JV\4-BD2]]R~dfy'^C{*D+VCZ}rU{soDm$'j+JBZa>l
    *j\BiXrKBAV2l{*R#a]*gqk_EjCvvTBk@?PG_olA>HEI3Va|mYE2uj&*]1#xTBeFdE?\u$XBo;Vs
    '5mmABw^p'l!XVrv>^j<ltovvBHo?{K_~$VT$=C1R!*z'Jx5CkYupTc-*[1I7;r)$G#!x=;^G;w3
    =YT=;N;EkWj'3>j-X5XvoK[>spv@_X}HgxDa][rU=w\H-p'Cw-G$a];>\k,|%I_Owxn+'G5>^}1?
    7vuV*EB*^pleA5-2zeK]X3YslVx5-\=*_RQ>C@7vupQ*JR;prn+p+BI{7WImQxH;?Qh^We?ERs{{
    G"KoTaY,RQ#1T*c>nJ[fpWZK_X*j+A-WVT]3v;>Gzr-ne2U^BB7rwYV]qepw;Ht^$IDXnj,U]iJX
    B=Xp'-slZj-8~'B~?sp=;o><_aQXQ3v]$5^EC7JBHC;~WAG5nE$WK<<5cf:GUKk-RVU$Y\$}xI^{
    z3@{AnlJU]u/?,!UpOIs\@YT7;EuiIm>il$uAO[+@a;HN=u$W~Xs]\ZnZTlBpZ^u2rEk2I1xuQJD
    zI?Y}x~J~_},O;OHTk5m'bjO[>*C{aGVGj(FZ'kQoH<w!ArZ]ei==V!Dl\$+cX\'@_{GwB/1rV1D
    <<\UX@C_C{{?w~~?^osY5]>5D3Q8VVkRwzn?D~ZzIJx5$nx7V!T<YzUwUe{~(K_=*j1}+:s5+]ij
    w]]WjX]-zWR<^*BmA[7OY@8VsXj=X\CVXU]>$CYz$TAFR3V?'jO{@*}sv!~o7Xp}I>j#kUIR@sOW
    ^*sJmI7YKsC+Jp'$kjeXS;[waBCG'lYnk\ea^7*K\IWXnFYH7H->ECR#zJl3l2qfz$8VXzY#5O7?
    n7OHr~an=kH/aD5xyrK7I1Im,j2~2BwKpuvv'WsO;V_kHw>pTV@\rx1p;~_OYpT,YX-lw-5?Y]^u
    vTR~-aXnV^pve!HsZVH_ii}[wKn[mUDD#w$D~Z+'EKH@>Q;L$3D>Czj!j2W_D[pa!,lE[XAO1{TJ
    *x$u)m[Z^=5[CY@*Ez1!>^,}2ox2BAnH2{qhTrpzDaTx'nKETE>{uaGBkeJsU*Q}#O*G@QE^,_si
    O[jpAV@Ivno<lmZa<VDk^a=z~o}r'VYvjTB*1A+?a>Vw$K\j&DDI1<jjzaDxoZY!'o7__hEW<TQD
    >BoHeZ*[!EDjeHkv*EUpXzV[@5^kQ<>l@3?9]mw-plYEOQ*#q0{>[Y~}xl-+,=$BlpIQJBi^*e=Z
    YsR%\_e^-D~j_$Qu;rTzj[$i'7{K{Hu]!{R>7*pZ7E{x;Y[{Y@rHY5}Z\]<ma]VieJ3XY{]WBQm}
    5K*m\1zeH<Vme~lK$xQwCER,DYBaB7^Ev,{ejQsCHzmV)5*15e]Txp-I_m]m*V1sX9KR-2!x'*BD
    213Yw*Ivp}"h@A[WBx{]mBn?K}T]O\<a]OQ@js22H*Ow5#;_1mI-co?<kYM=>m*r\DV\<}^kz57!
    _U[Doi3VVjOz,Y}m5ZE\XK-V1WAvwK}B_R^{,H5[[,_i<=?!=l2j<w!yeC$x+]k2Z+_JiEe*HV{X
    E^27~}3CjeB[*=xQ'HBK]I\,}?G-BQW1G'Gz2RH]7!m1Ovje*Wa}IVVVsYRH1GY!Eso+CY[^e-D1
    ZGn5VsYp5_1@I,eAv2uAgqu]2TtB?'ZrI^iqC&^+={$=#$nnJjU5Vji-VE?{;[~UIn>o=E4"j]5k
    B@WuKX5OVBm^hXOp}{Q@KGi>=$;EJJ_Hw:*{5W1T7'V5>}*Ts+o3Xol>[xzas=u|<V*wxI}GZ-@C
    s+J@V<7[W-*>i1C#IpjA^,!T^BsmU_XA~o2~J\G5$>GsDiEZv,w3vWDIx}'R52=$~vIJJB_^]ID;
    VZJTRUoZxC{-\p{X^V#1Js#TGA$]TwsE_^;oAY!W[@E!I^!x_To{Dxm'Y*vE2x~Oe_HpbE+jnRX\
    vpG]7plr5v>1{<DAZ53v7Up<?o~A~CQr3E3u,HBHnBT7wB=#Q915GeC]#T6,Qse[nIOpro5xEw?r
    $ECvAu7Ep>>nl_QW7*>v=-H7I!]%7AYmxp}T4rZTem_IE|5EwCJa-r\5[KxA|B;-CIoiuiHJB[Ta
    ;$^oRAU_3vYPO>ORDZ;Zp1T~Ez+jO2ZO^=v\er=XsEx]e<vw7m<J>_O[mr1oR,K?'X+ep!,Z2Au<
    %&rXQk2Xp$j}3!eb]@+?8i=J7CGzs,srsF[RU_3aoAeon~.V$]@x=_JL1*u]_el<w+z?pTAl]\e-
    K<<IAC]R:koYXRm>+w_K'}p[a7Dnl1n1!G@l^Gz^?NqpH>,inY]1;{]kQ'zzY@?BlRp5@nuTz+7\
    wEwe?XBGRn7?p$!pCriN^$$VKU3zH'C!U<=#ARG\AC=5z\v5V+CZP'eI'*>G;_?^Z\Jl}=lj}T\I
    ,,I^_~HsV<-@u?,w'pEr_S,ZxiPQ!-WV@B]}DewH->_^$E[DWUvCuDr'{w@ZY^#*elpknBT55jD_
    }ArsTK5ueR{:sxv_<zH?~GDK,oCW7A5?3G^17==>@Oz^V>sONdW_R;PYHnx{]ZuZA=J7nHD3sxV^
    EY\F357]jewz@GV-2$B<\z>R5U='+aGE~B~EU<*OIR$ayY^r-L'i{@cz>rC-x{}AxQYL]T7*!Q5J
    RLAoe3Se]Ik^AnpQX@-x@*@|]DBoiBej}#2\;QmI0V!ve^5a,$nRUmVB2rE7\pk>3j#\RHpUG.Y?
    +m%v5QQZ[AXyJa1-5O<z]VUEZzKnaR^,u-X,1-AQreXX@DriH_3C+7=-rAC+EaxiHBY_p}asDxVR
    xjE@~A's,752x31]Y}'?CA_1q)lOAp2\^-p]J15=j'<S^V)v1DCQ^op5YvHnHD_$\^@II3EIG]w=
    {^$12,@fiv!}PE,2Z^!EQrVQ$YYp$]eHl\[K'U=7<up]WWTuEKY1QBV#Q!{]iDu'[/JI>IMz2@\o
    |'V!*J^V$a=$3uD!GiV!T}A+3=QQDmwRkvsDOC^_$zBoK6ZauWHo]}VDH3EI=]"G-;^$e[Va>mKU
    7E?s#AVzeQ^v]VzI'O;C+;U9zwOK:a=\AIe\Cw73pM2p>W+_2pu}+Hzk$OsD#?$B$C]Z2\DYaB$H
    JK~=wn2oW*?j-EkTJmWCA$$B>Y!C-_r^p,'$Dkz5AIsj*'~.F.DEsa5$~rRWrW?H7^vKe>oR,{sj
    >JeGx1/}x#DuYv<e_A1m]$kRL$1->NH[sG]J{;{*'$1R{1pHu$a[WjEEBeKUj@'}xnvJ_r}XnVwp
    Tw=UuazVC*z#}7lkJ@H{,>x[*{*7!D,_xDF{B~X=r#a^$+s~$I\fgl_TxsxrwaEI,3suBI<]p:+T
    O+1>J37G+_HY\;?\KI*e]wIJ5H7ER#>5Q3%'R;eApsOVmj[1ZA~f?vsR~EU@2Imv]QlRxEWQ3l_k
    @aUK\C3lC#O\FyBz>'^AE]y7$1@Z-mA-}@DZl}s<'DmJ13?~GuI_2VXkVoYvum7,>r1qtRI5a@+r
    z]p3A}53]G#|hjo-v]ABZ
`endprotected
//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin
`protected

    MTI!#@v?m#wwoWp{aj\Y=*U[rv@$m2'\~5Uu>FLQ@$[LoxsoW5x,g'\A@[O}Tok$Cej*Y3=kuD+A
    E2T-#vHARvjk}]irz!w$wIi@DFzx^QI}VCX$sD72[l|W'#Zz1i,F|,*Eka1#>Y]k}vX}BJDQ2-a<
    ]*QK!WIs3HjC}75A+?<7~H1+pGuxsx#<B:[CZ#K71mD7*[2jluOB<<*E]=&}XI<Iu\$$m=_?1G<v
    a2CmrY?TRa71oz2(vm@@Ko*_Z<AXZ{r3UD+QxJX$_{XzTEGp#B#3uC;V3lp{J$-[!a-QC2a3U=r=
    7wE5S$T]EfsIX$rjl\ea>e7jA7hU]Sp_3VG=*EGT<j,ODBpwp3i|Zn}u=~W'@ABprzEVbK*m36}e
    ]_^#z><Ix$oxw,VH5=sExw?XGux._YaV%^B1m<D,@*EVrh*W_V{XT:,p*1(}C*K[eHaOKz5$W>B-
    C~zG[JskO*7o3!}GsX>5sV@;D~'V=A-gDmZ{izV-nCZ[G>V$;7D[KnAlF(O#GJkY~J'>71)z51[J
    [@*z$_Q|hNI73TDx{=**O;ZUs$-^;,JB57nTQr,;2Qn^HA+>wkDmz7d<>v\kB{mJ,m@hUwj-RA-R
    KwlQIN)?YUZ8#[Rp{w~ar]Os,Ri;}~l+^lV*E#[TC7!^%fI-1WomaVG#\lB+1k]RYj>w3,s;r]he
    g$=mBtNppxnq{U7;^T<{3Yx='[?B^@xKz]?VGp_lskQno#z7<[<wOgJAQ~T{,G<7E2@Y_1bG'irt
    jisamYk~}BGD!Cs^?TGZ:[~!kAXoX^a]xE^Qo$WU_So_BGnU^=wXw?Cu@XOxO^5J\ZBmW+jW]^9(
    ].vC@o?EiEiszHDD_[jn1#_en'^,TUEDCG@U}2l5[UIGjn\X-3geYQGvCpk<}e{2]KBv]@V+5u\[
    32aiVEi5kTZ\,xBeTGH5DG27=p<IHR$_uC=pC~,YD!?IZ${C7K[==H1Q]Ce'v5-zx,Yx#5=K1wV\
    u2OiX;Q*;A,ZsmDxBk#XE!X=IiR@aj<3=HBirz'#<Ze]5pv*XrK}VU]lOJUrp_pCJKZ,2K[I]e27
    T>;3];\0['d,<11kHVr]j*AR!x^tZ'R=4VAw]5w>VZOn1V35@Ur+-7W'=<+,1na@n\j126}!-71Z
    [;}JTZCio=gYgp3}p2rQarWaKg$%Skwz_UzOUq=K$JJDre^o-n_X@s9vs#ox&_]H-BIU-~{>}<^k
    };<n;mH{um1KW$+Du8#{Ow=/r=rABy0jK}a,UT<aOzlI<mQ<rAz_KHYRURwcYs1K7XX\x1-U1o<~
    8Qke2?[,lJC=YKsk'ADpIeBoDkIO>C{eK!Aj+Y\]HV{mj=YBIm$_*z!Ujm*EVari[ir#![[]X{}?
    ~XDp]YCuW]Q@eG;{znl$j"%[~jeATBxp}D}lZ{@PJO$ERrQ[ZRZ}s*k-=^]![noEsr{m]z+!7b5Z
    ~aTD;ops;R15*2*G>-$H]u@[QxxK'ZQJl'ok!B{Bn$>wswXG,-W]O@E3-7rBXoK-7DGxr{l-T{{D
    W=L~D=K}zrE>E}^A+[?V=${ZO2U[Vkn9BKDp1xGvCu[RnY-1n<es@}DaK7!;>Go<L3'>em$'pHC+
    r\#K,cOs>?;U;+<$"}OTX$e@U{5T=8{Ba'},'VnTnr][']UU>5,?+rV'QJZ_vB>CJoJO1oss=o8I
    1KJHC#?$HTCRvev*O}p]2sBH'ow~-1jlr;YR;\+^-z*D?6{1@T-\$'tz<Z>OsBs']wm]i}B^EpCC
    ma!$-OJ-\3]l$D!Iwuvp+ssZ+$[taxeQ~][!Ooauj<J['KR1NmEoR{<erH'ZZ-{R\CDKOBJvm,,k
    3]VGVu^XGe^?GzXXzrj>*JYme^H-nsB,lxZn?3DVlW[}*YJzKnapl#T_E^jzar+rr~I{>/HlY]r2
    ps?R\x?'kJ\tKwG=$u'JGJOELyg]zOVB\u!3T]\[^u?\#DzB<-[{}Ez-DD7x*#D}n_x~jT,$eXjI
    <x<'l-*'T7]qs=<!<wDWxC?wpH<D1",U!HZ5GAC;WZwQ[m}%ajI]kDnrUVApPc*G7*yYGT?;]?B#
    ={IM_?lijQ#Dv2VEH{O7Rk3eq[lz]N8^{,IHaK{*,Hu1z!WfSm'}x=ZX@BJ'Rew5k++G~Y=*VsGe
    i?5+A(!\}3qGz^T$Qx>3HE1TrD#ExmHixVYJ[2I{ETAi,7K]+p\GkDAvJrnwa2YC$_uMn+TUkDx]
    ^RC>eX2l$G}]z@Te'zUzjZ2pT,5Ga}*w~Y}[1EXA\IRvw[H,~vZuXr_3]X7*U\V-lmlBDATIp3a+
    3rsErG;vz}RlB3\KAYK+u^'Z>*$kZo^\O*5;'_!wE'j<Jx$3&^OQDv#;nInO1s,~DY~^2y#-x;N$
    n\X]H\Al!eJ]5}mKYHAQ+_$w+A?i,xHK}!\\=[VC5E$G_XKjG$E1i*wlQn{pw!<yov[7k>[nKGG=
    rsjV2a-Jenu-*s,V'e2@8~'-]!,A{Q~X\oU_!@B]'seHxI-2Y!r-GTD+eojXEmEZ\jsa[BoR;Wa<
    Ae!wTe;Q=n<KJ'<s?i$rr{enInnl5'i_JCX*+2a^V@zJxADKKb$*nCQ;Dp[X7J1+GY:D'5>IW<_m
    B]Jf=m@Z*OvCC,}5a>2x-V?@m5$W-,IAh>s{s%}HBzv{Zl![}i[iXYmQr2Q>ws=$xa=[1@QjHkas
    n8rY!,lgjRp{i$~#}xk{75XTIK{wQGZBrp>]';IZ+UQJ}R!\X]HCJ>C>a]jrQ!['J1#WV!7O3Glx
    K_Yv[l!{'#1>YYQZ7b{XH]E>@]A'2p$EiI0waR-$5~rBA<*RHJpyepsxHR!?3+5zI?*a3=Yl]XGs
    xeskU\VK[_}j]\Qv1RkB)5-]RX\EnYD3'eAm,$--xK<CujsBzCVYDR1Y,dUx-!t_Apl^o~E7pApn
    XQBm7Zl#,;ks-!<H,UpYpis[s1,_GHVkO@VHp?DUB]rD?9G*rp_@wn^K@Z2v}v#]xJIAO={V,G\+
    C72j#B\*_vCH>Xvp$J1'oVw+,A^AH?'Vv-se3eW,R-]Dxo]QoInn3rjTIj1HXT|ksI5$-KXqE#!?
    _$Ce\mVeVwQ3]7}E{';CJt$1wQ/<GDV<\D_oEY\s_>WzUO#[G;Ho\>=pBJ$C_^p>],v^{1YDX~aw
    ]Xjmj'}zoJGOAKa<$n$5$GmWRzVH+C?''Y#H'ECD}B[*3lp}GTzPlD]TQo!K5#RT3BU@hv!EJszB
    kU[X<7~UBCHE=_sDzKjwA5{rXpkp~#]\#wXem0DHXw@[<^HO{s95JY,#aQ$Z>Vs_7rXXI[nBrw]=
    rCZv#15rCB\D@!eVMG@~QI1v{fdT12nOs<,7=Ip{QYk@]<[v<wAR~lH{A^Ik5#]Qf-GkIsn]IIj+
    __H-ZRR*C'ycA[a''DVJ4kEO#8]x?$xs*Y)=FX<*T\'?29>zp'7uK^^+,s1>\#\71]n-vsG[7=JR
    <~$Tp?|EK'lu{uEB3GEnXTkm}ZT\C[W#7*uI,A@$Tm'Nr{-DE@__]G'RnlI-373Oi]WRE-$K3-~w
    =DB+kQI-\k!>rR{~i$}-mBjUeVrjaD+O@U^^2^++rl5W_<CW\C*?k<>!jYp{Qo#Jr{lnn+{3Cz#n
    W_u1T<;Q7Q_]U1\xtn_R2reK}wECliY~o1<XkG<XV}kD-$*VxvT+C{z5$UDK!/;VVGs-[}\ovCKX
    _'F'n^_V3JICb1naHz_!'7{YsRo-]upU[k7>;Ir;7o_?nxnzHg>>$kBVR#?p^x#vD=1{{=X}DecQ
    }H*VGnXNUx*kqwwxwlQ5Dww{'X_Y;bAYsOwBWKw}I0Us7{ZD{u$z+Kjv\$?[Jlzr>Zo+D]5VviEm
    r]wjYpp[jX(aX2DslIYB#'_uaB{-5r+[k'=>n7?|;,ka1$Exl^kG$Pz\xHzw,^.h@-QeYuZ#k[*E
    sr)0QD1z?TzQBxuRAQVmf^$]#NKwV?qW'pp;}e>sI'B}I^n$JQlmYmv=e-GGs=u=TrC1v'wJ{XmT
    _w,jk@U=xC1@Ba$D\?BaCY1Hl2+~ao}.Aek~}$UCo~I[,Qkj#UvlxvnCe>[>?<l[=K<[p*n5#Dr[
    }!,}Up;UY'e\;Qz#\pi!]7X7pYHj%@$H2OA'[G<U{]#!un{]<p3~{GuJuoKI[==3A}W-xTBI'pD<
    ,Im7$Gno^ooZ-sKD![o+z1]e}3UQU;<OO*VCT5>nv2=^w$O!X3I!oS,@DOzs^oa7'H1;$i}G!3v#
    +s;XDJk[w#6kx{vBi!2C~^x]]I$sx2Em*!1\a=mxmoiu7Q$A5Wk3z1EL<<j]O\OO;>AD$pHobO~Q
    ^MUrD~mxG?;*zr3,TxZH~?'2{Gf#E~rmCkxdcjao7z]O[@G=Ov$<UV]J~IIEsn_TRtR$eZnAzVmR
    a]cKUo,AO@IIWD=2r$!r$\HY+C[_E-*i$~Jz;R!nG]>,5^=#Y;$'--#8@OEJ!p,Ul]]l++YCKl--
    *E-v8pio;W_k^?[RQKQ$x{vm-,A<+U'v$\i{R!}>!me3vTV-@UB2z?BA;nv~Rp{{^Enwo-pa-$Ae
    !^OGVK^usi'$}G?@-D[[l'zV<hY^aH,u+J@x?;glCB;-H\I!eYR-BE*'_rn0Ha3x''T^zGs+W='A
    [1ZBR1mu;Yu5?G;=rTRa1#u'{\A1Im,ej}ep5ejj~B*^OWI7R^esGII;IpV#x+Z=U,3k[rE?sX_i
    yQ}*_C]?{pvmQBWeX.uvK,zK[aQn'<m7]oTGl'zJs,!XB7mw\U^C\J*CRs}Co{zVu=!_AWqGTElr
    BCXwTsY^?!1?oIvJpZ^vJoGG*-EGp3ADBQsWCp5UwnYLL-V5oX5aHm*7<pn2A'O<YMCBCV>$[5Yp
    *Dh,~Aa2j^G3e~+2<KQvu]UPe;Glp3u#]eJw6XII7eE5OD-sU,7>2[Sq2Rz=AI<ur,*'V>Y=RfCG
    3aU-[XJ_JZ%IJ,'cYBiRZI![5JI~TYAQB7XO*+n[z#nC{\>l\7
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#[!rOsannREBOVWsrh^1CUWeQsjC\>E__[V?O*=~o<s'#+[;w?#,IU'\-w=8nYz=l_;XeD;m
    xQK;dX[+2U{){Ck;G$k\s{ErsSKwJUz^;};<VnzxCXX{DwoYa=@vvpQR<>lsW7R_,#5JxC7U>V\$
    kG*+E{8lR~zl#lEy,U^@k<o~BXB]n<j-[*EZ-YDvrT,i3-szUOAn\!mw;9'!Z<275rEs;[OI;]Xv
    R[^BQJ][{Y~{x;'3l3oi+#{ouOO-H2-r7B9\HY!}lk]zE?+n[<]wwn]}^31}!I!*\mvZVr-Tow2C
    !>mW[OvXwJKQ~->>XJ[^AAU1$]k|-wpijN/z<_D}Yzi5i[*FAn*@(+=wlN^*2<^ZpV,}<<NVO&X7
    ,Jv~u+?[peIK*2:o-[[as!Z_>m2Y8;=#U~U2}!sC-QinwYi^?|_-@3a**?fi1TuB3Vu5B*#;xjBQ
    jes*GGr,Y*_'sz[opXkwl>n'o=as!$iY#3\Bxn$o=]2=OQopa$1pk;3#C][,R=}@>aoaoC^H=@+{
    ]R@skUTH]Ga[6>AYG._VD,Qzm=>jUBZ-lAB,rUEvo;vs]u#H*Tr#Qvl!VOO_<2DIn<p,'e*#5Eq!
    HZkz^-w_s$eiYOXG#UpE&77kZGGvVjX*jdDrA!+z+n3__+UCm3}OYX;[lk5_<A#_u;@$!!?}TBvB
    T_GCv*->ACzf2o5r*D3$Z<W},Q-WQL<<53Jx!<-IW=37@=lfBJ{=aAOjW<JT=@X5c1v#?kw@;sAK
    wvQ-]Qw}\l>X57IDH[?'u_~BQ]]-nYHWC<IEp~BC!S<=xY[r5<n7u=1;n}@=ls^UI_!Ic!zH~r\5
    zW[^kj5YAU{vAc{]@ZWp*BBH_WDaJl3NCQA77BQrv^ArPy&gVZK@,;DX1'vesJKstOKK\_vJ'Do\
    _5B-[U}5\!'2Z7oW!;[l\\oY*AIRIET_7p{leyHD_GkU5_uX_1LZ<ZK{B4x>WWX$s#YpAvxH~_X$
    @W($rZ7G^io,Q@\[UGB2vW]>UC@RIZ+G1^1=V$}Y!2{TzI3}a_^}<ATY]Y{p1W@nx{Kv_$!<[~l-
    }iG5]jU$$mYNWsQ2Q+O<7UDY,J7z~1l]e!eojk}Zu}3B*1Az<Ap{crZ}}ieY*eV8pnUu\*VHDGj!
    p*R\UxE=ir~p/1C$Jq[Q\a1aovM*QoCw(spjQm1D-^]CxA]{l!z5@jUa<T'EJT7oj~E_Rs?_i-r7
    $BI^Efj!TOE='w1i>R3}ulk+prY+Y-7#QRCis>+eZu$*3-|0{BJ}i]?l3^?ophI~XBlTB3f,5C}i
    Cuj9QG]]~H2CZ}3@r@TE<TK+e$=~'*Z@7KIW>}jVsxu57GkTaroA~]x'CU]uD;-suG;$x!]s*Y\U
    ,~vw^;KGD=,u+wxUOV*{5\lTne-VoR*\joK@_H=}ujWU=N.j}D=[Z}~EWY5$!7vBCB7E,#W?_2Xv
    QGK?DRBtn*U]x@^<kAIa,=]T{X{rvv<Ze#En3s?>u>7<1w@TmoYK;B{eDmW;'Upa!Hjv<|rC+?B>
    G>R+msAHZ1.ErDDAps}p?\1oj\!TED~Kp5=-5C,=T<!{,'V|+xppUjBlo?A_0C+rYIuX!5_]K|En
    ]![C$zUrTpHC{E2s7ozB^}ejUQ=D-uT<}o}2<3)|{}W[<wp}C#D!XYiY+T\2s?KY2z77s?-VuC=i
    $A*I~]jVB7TjQERE['=nA=^>p=O}e;o}s?ORuDQ'XTYmAB;\*;EQq=$kE211+YJo}OxtB[Ka@C7@
    *s$'D;l?Q@72Ey-n\lQawp!Xl}2j2vuw7QRmVs2I[>OHx-Y-X{B?[*'I]mQU*-{[QVVRA{f@1eXn
    aeaB_@>8;oun^W;*\Y}mle=Jl<u2l^EkiII5^E#K_']Jx--_e'j2&T+WPknm?{Te^e<!aWUz?3CJ
    TF=r[,:7,Gk'J}\}w-$m5V{EETkS.7;ra}(kxU^ko@_'eXx-5^H7HQI\<]T}iaHoHHj<slItvRD$
    GCA!7wr_K5,*v7}=@[+>$/>X[=Eiva>A$U7[{Gn}Hm^oW!yU,Z@Qr5V*aa\T_j<1BenX]z#K$Tes
    T+K2n*iD^z1KwIITGw!6B,$7RGu[7#1KBxTHQHj-xzz@dojjCp?K7}_+U1lo[p!;T][GHT<n~s7~
    !-}1-]CT?;aG_PT<GZ(rWjOzDviA7e3\Q<@X==$~aD15EC@HX@;~>R_'WwnLX51TcT5#^?Czp]@'
    Q6~xK1v{lA27x5%G<[];]i-\$zi*]J]FDmoGFX\$zQH}eR<K~>ox^W+w'%)~$a{j\1[a=eD$^s}o
    E@R'aulz?w,'^~Z7G^n]@vu>I3D~*X@3C=O5[i[C+}']_BH-vraIIRZQA+wo2!JXTI_KA2E8|-Hr
    @:HwX\}QVQnV-Z!ex?Z]?ROY}U7Vr*m\?wt2$oUWBv'4GanjBJEO$V5=D^JA*'zH(UwO27rQl#r_
    _\aIGv+C?xLqe5sAHVQOU^A^^\]DnoX*v<e',QZ}nn~TW>+13Q,Wb1J*V7!{3<<j'7E}s_iEm#e\
    J}}B}/[W@nm'1R{Gu}UU@T[;T13,'r!$[s$T[v1W-}B}@=B}'!r'~si>^$i^zlJ7^Zuz#Gez$r3H
    mkW[O!x;>{p=jU\5A]W}wawD}r:d;ATEJ-rv,c+TAHIQKY|}JJWe=swnIV'vs]D}G^;*7,;'Q#pQ
    1RT1OV3=T1*\+zR\;Jp{7#~B@lua1?UX'O<zIKsmxo>X_?7DaX5gHIU^7Gz+HD_k+H@pO}+-X,]U
    x[i!z<U@GiG@vn\*B'l;vk{n$aCWN[b1l;Vkr]C,j~pl27w>>~@YkwJx3CuvO@XoCp3I;J~'3\<I
    HwOz;BDpDQ,}33]s^re,ewokUp=?_5oy*#2J5o\{3}Q~5#e7QI~B!+*H}ezulj$2vpwn?[=o{7J$
    3jep*iu^QrUXxuQW2$-El5X_+Yi!@[j5)[I#_?=E$VmCGOz2?G!D\1<u*$k[_m*IK<>e3=DnV$>E
    <Un\{H>Y\jRn@5O,wEHuzKUo_3$I$m7hj?Yuv!=HC{Ra?'{smXV!xH+Z3'zmRYQI!EHX~7z3s@7<
    ]B;GG=AvR*#V==\o_nZ@bDomG1<XOCv7u{}vo]$5ll$*,6VX,AvlR*\ow}CX'll+=Ti$?uI;V$G<
    j2ypwe'er[<sB$xLnTQrJ-2,6CYJmxrEXA=kzBKA'$~^x~ax\[+^^^X;1+Q;~bEH13,H~,,$TVx/
    $<R~=Y{Tko@vK}'T0#TQKEY_UpUe}^m\V+=+Ge$R2C6CGRnpxmY0<,a}[izT^iGXEX+_zHE?1pO]
    )hi^Qi*1j_]2uR<s2=T*1;+YwaIA=TSeksQT_?Xl,_*GCG,2*p,^-A;+ER7^]p7?,Q}JY3;pD,B5
    oQ*35}v5]+j<7m@Bn}pQlT*$<$kz\1pWETU,O{E8|$33ERxO#p\;,o!^_JXvzl}IjkVAC=xnmQ3$
    [^GGKj!\='JVKDVC[RIC1gU^rj0'\]i/%EGpaaaJ_\o_unGrp[R*mD*xi/DkEknVKQ]uWzrB$EeY
    {AgrB3#\uA*;,AEs>OI<sWkv<]~o,'{:kv3@#C5$J-{-J+m>A_CmZrGAI3Cl__Ja+A;k|ED<~[,i
    O=~^_IH\-sOV3XI{HYB@~pesx}?mkK^lmLQW_ssxi<1sC~Oj{l/LkT77p[RKrTUlr$3[k^B5b^in
    eil*=oH@sfmxHs^5^s12p3BrO^*5EuBz#axrW5}D>\7'A<kVD;O,5ev7_A0@D[p+5Rpn}Z!plB@=
    \?H![}?KVaZllRE]OjUlR?;]llYC2E=6-E#ll6I>w1XQ2@lm@IVlk^ApOODX-!TR,@[F=WzmBpJ]
    2<}~BeZKTj<I1<7?z7?JX}{A*8rp\!a}v-ZY@Hs?BowrsWpj^V[]I]:BKnB-Yrl^@pCi+I3*n!W?
    IuZWElxZIaxOEDE4,R3!ll_ix3U=RY!r|LTR,ekO\$epRD"HxW_C@Wz5lJpR-j@GYCCZaQC5F3x+
    Wua2~SEYO*1=1=}!;}m^Op*'^[cpW5!r'ueZVjw$d6}gF@o+e5aHn[emI]oWrO3I_7^-}K<[Yp$!
    nUC{V1HZ7OrCm>z7@j!!7rkeskD5_{x^ufe-x!pu<\;v'{f5rTlCmwp?<ekTxQz]Dwz$*a@>pl,e
    YTE=plu~A2<G{;A='}p-},$G]3>eRDk.*u>svv'vl#~E?s*U1?+!Dt*o1VKVr;Q_;Gfz5sZ@<Y-%
    gHo#K^X_xD]aEDp[}<-ru'$E+T7x{}]ZAZDHCk'Z\j[Qal;IDoe\$,BXjHEYJvA}@$tOXGJpT2l1
    W-aW1}x#T7'sx'Hj=ku^_YGBQY@T[ll#1Jo<awnv\ABrROuXVwnlT4)YOHjw7D^G[r~<5AVH-x}F
    -]+ZuH=-{=IW2Bx!Y5vkCQzJO!@7@DrU4=1jsEXQv-]>'DWE[2YB#Y+-sD_7{b$DV'?ORDx}G'T\
    ~u2^YTqY]E-_=B~2}l>E#2m$Km-|r=J=R}GsvaT1uVn!R[=^%,rA!6[7Er-[7A>*se:WwZ,rz;>e
    GZ=XB,-0=\e$^?p~$B[elA!u1mTQI@<K$QY;AovRh@RA3@nuE%kXDuro7xv2-<G5<_D[_^\C?\l{
    Q?D=\D?'G,#X<5!}-o4a}l71j[31${}-{p[YY!sD[EDv-@VL{5R+]lUuR~-H05J'J=-]}czmp+Ql
    D-lf^u-Q1-J?e<2#I}}Tl75D=-\$x{,{Ka37j5Hl>^5DTD@{2e;>aj;WZz+O4G!m$vzrREAWJIIs
    ;'>QnrmO,TG1!3a*HG=Cri-z<xiOu'uvDwR_O'X2G5sQ-BDw_@^;$BmomR-l!B<neY-B3n^\T~VD
    $J]nH,Y@Gbb]uQ@HC'AHo@ae;p[wE<zwxKIC5a7^R_ASeX;B~=*{ms{GEO!KQQ]<qoa@'],zj\Z$
    TT=v\]\u_IamQDEG!^D>mXr-ITE{RoY~v#R\$uG$CwUXJ^;ZxHpr2;E7Ilv;{IauR7kHG^jjDH=<
    X]V$_SI\o!a7@-A,VaRWA-,C>\3wQ]Uws}D]}~op{YHj@za}3[+1[j3+wuu*<ViBpZioYCYWr^j7
    K,0"^s}wj_278[<Rm!5m{'>^$*G*]}*=D21Y<V2A1+^Er_JlWpWv$Aa{~|H}<7nU-U5rAH^n-u\T
    !QYJpw=m7X6r@$E3I*?z2joHe<1R3D5|Q'#{rjJGtKQEenIeH]w^p*oo;fn^325Q<2H-}~wQXR=U
    ;oBCEWwDrK*Ko+kCxB!z1zO+XUJC5XE@<DO'7^YOJ$Y_i@a$uWpXT\E?@J:+[OvE<lI#Ur[e~Vwe
    (#rzJ>w$?%Un;AeB?s:*HY[132-,X'T-<![HY5;xx~3Ri>pAG@~k'O_;j\$l1pnrTj~Be\>CQVVa
    57T-r<^OYRzkV@1aXO}_CpYk1'$)gp+p]~Ck>@E;VYk_!U[UX_*!l2OAvB]>^xsvE?{nCZ1#;wsA
    xx#G#5>U][aanOI{Ox<zuOW~wG7,J5O,?$BLiXCwR[onR?Dvx<;JX[3rx\aT~+2]Te]pUpA^z1Ga
    sxDvwA$w>9<p!k,K>_Z<!UBK=D#vskv$e@RWKsUQ#{&c\;r[?=UO2-=A*w{p\l5jz0mwW,waQw@r
    UXx~;E!]?!jI]!OBu!JI+p1Hm#@OoAT5XowH1V\z5pVkDuJ[r2^{JH]GGRy"-7xD61]Ewh=^w}fC
    ?}l[o]-<'~UsnR-xr,\\3n#aIja$E!2e{Qs~pxXYrZAvlwD!vIzW,#kK[72Y<G~>v+VP#s5i|D1Z
    eWx{?2Q>w+r}=$1QZMCwTlU]n##-lTZv!OD+G*55!HpDA{WeUw}u-}BZoT}Z$Z$rpoq>_QaRz#}e
    mnxl2T?%rDCX;l3\jpp,B_D~7>,2\+~=,_x+,J>DeR,1]3_up3l7TC\[2ejWBQACd+}a$sXHKT(!
    _e$ox@~pv^E11{jI_@@fkYOH,a3p1''$AD-p1?s>zJ73zBD\|*TY>&O^>jD+>IQV\Oom;J^>TW@B
    ;zGRIQBa;B8e'Q>E3T?=-=3^Y#'~+R*e+BVKQY~$VAe=+EKOJI#VWv'$eEZfRe7\3V\s~$xis3}J
    aQ7J]'s\~{J*z^WIj@I@R'1jA<E]TTeZ7RIr\AQIA1mYI}U,v-~u3<_]H]Yn<vrU*(BYHX}v}3jT
    \EV%ap>z7_Kv8!1oz}3I-:$~DwQQ@U=*A2}x$~E-jH]*_eC?wui-*TvTvB?}sk#^ECeBeAqPtoYR
    YJp72Y;3ZTBwX$-!-b1=~axO$#';EQ,Z@^'#1]9i-=>pH>C+Iw]#>R*=@Vu@$Ep=Zl-yDzT]g)KC
    ]CVJr{izp#-wU2^SO;j[1}!Z[i
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#l7pOYC}_1W<lVWlv^gs[<+kT@wXYr3L"[cA]i}iod;Rj>!,2!w*Kr<5!<XY,=l_3XVD2mQQ
    nO:X<+2U{){Ck;G$k\s{ErsSKwJUz^;};<Vnzx#XXY*-oYi=a<pv[,7=-rka<jwB1G!>^wl5v5k'
    ~=a<hWsmA'Z>+|\U+olD;r;soz=<W[J_Dazlu]A}2Up{oZU7in~DXC$}@X}],z~'w$Cf59=CG*s]
    <^<nB{HCA-T[+}^\EBm[?*n,WnG~C1Y[D=#VbA--T|-wDD[uWXQG*m5+z[zQGB[z3!fu[?$BIxUo
    uj\)O3DvuH<IL^U[{;7#}Y7~-=pE$CGriHT^Bl}[O7YvA^X,=^3pAk<rGR\>BD~},Cu2eB.6Ek+_
    '$QO]IBol5~,g/>pAG;\TOVTw}xBkKwR!=fNS$F}mondY5IUQ^$n=^,ivaT,Gk_#zs,Rzsi!\lW]
    I{C*m,O{,$>]eTHmW7eYCxxT?,YpV=#E0GzuZ=~v[-_zu+DA~O#R]lzYnRD3'2G=TE^B#Nk7V]"H
    5=laYl35Om+uDnuEl?s@rokl<@=MBu+KU<Q31DxVNIWZBio<YH$z]=mI[97vi]?}OT[l{e;G<CS|
    ^?v<uGu3=D->Qn[wh,wZ?;U5WzkoTsV[maAYXIdIQ'DVxAv07{'IBe=;voAAB+oEAHVU]CB3O,G>
    =e[{<*lZu=mufV3;nws[Ie,z3IwX-I]'Iaj<\rK$v+B>sp=7=Xn5BrE5TJ}lOnw;A+1>=xi7{gxr
    1JZ_A-BW~>H$UE2V#G'W-e8oSx!+]O;WIRm{B;j[~rKZ[rvT?^-R{Uj_XITjCaE;uhJsO}E2;,la
    'v}{s}='1CL\[5#c#zG*mUx{{U3@Fn{VCR[TO&Q8Np3vO_,E37-*\v{~B_w=jr\Q+B?p_^g7o^Q}
    !TA$CR}-He@VV,D'lv=!1?kK\IA^HjJI>Ou$I^a'2X~S[y>'G;!=1U7$~oQusDn{!mBLn7!Z1@~e
    %fV_;us@Ysj+2mdzG\w3-=!5'KW3H2kDpzR*n2nV*Zezp@u3I~[v?T'et^^jCwB[<ZziJe9xJIvx
    aG>zADx;6]3+]@vHw!sp7QY=$_m!W=zk\[A_@,~@vQDK5ovJjk'W-T^WKGU+)p#;zr$[D9C2TRQz
    s{cw'#X'H@o=#@T1G+]xInnDQI~1r{AjX{wiV!UB_uz471v2Z[]eBOjU't|+1C@B1\;]zXmz<_#I
    1I7t,RGaok5^emo7obPzwr~YG$+,U[_ivjlr53^9oCz@],UnkE*xn^WOU}<W*2VUD_jm!\kZskep
    tviu>1H$-_nU<[oW;\>wAu_zOI@BD8737W=5^7Ie117O[kj]'~RB}7IDJ1lA*UjE^v3,E;rYJ~w\
    DAnjlo=o{UHU*H=[n,jX-^CQ!vj3,,KDj<Ye!E]$J$JQ,u?H}1_D!_ZX_QiwnsL1B\r:ATm$VWU[
    n[Yk7]3vGC{oy,@Zz-HWB\s-Qv<G,*GDjz#Ra^@j'{s};^+GXQ,=+*p@xXQwj'BQvQeDJTIvA5#+
    *:bnwjn{E*o>-TT]6pn<$WoGZmD$Jfu>QG@1E~5~5TRiCZLWA+\G$TJBj'\#[EVz+$nnAG7GmEnc
    G7@oVmNkXW=?wEBl'zk+C<!J}YXkT7!<B\!)4xHl-~z}ps?2E-=V-@RkRCu5KQIE[4Qkw~JRz1/"
    uaHI,el3?RiBNIpKGvnu+!nZ}$}pj>wp>5<}ECI*QO3IjQD2nCne3!D@X&$a_j3r^Ql_Oz}Cl!:;
    pEVa1wU[zYCe<D'm5#siD@aK*iYb[mr2G52;XQUlliJDR<\B}BKx:M{1QK!>A^z3IZwQROv-w[rp
    1aBD'WuE!T&uHD;MzEB$zm<A,3}+6W[;?xKQHS$\$J7+Wv^#}-=un7#+Kr*KExUB[=e,Wkskj7,%
    f.[nmB5\^2'^iEN<A5T]vn3mXO<R3V!G+G'I-H,,uOU]CWr[ErEloH>)|Q~1*)m}7u:]BN;v$k?C
    ><pv<ABev-'HKxu>Yn{BV>TD=s=*3nv$WB?z}!Yas,op@jI;RZp3D[(C]~orrE!wX{O!{U!wGi>3
    zAQcU-K~#TK!Q',!H+]$xD7w']^;zwD$*A5Cn[wB!TTBQ$zXC!)7XB157*29#CE=G.z$Y7I5>~*R
    X7lYG^,QKvMo['^2R$T!U{'friOQP;wnDr=5sJU+'ZHP3px,F];{!^&XC'E++AxW8-Q]i!RGr5v1
    $I]2\>Um]l$TpD$lwIO@}PJ]Qe&Rk@{-\ou5UJCA^uT[2El=w-TOBEr-UX{!jvmODkCD7-o@{rsQ
    'H*_?OIk[!QV*!k}rR@ZDe]I$GxjGOZ3152*tX7i}weB=YC$7z_kuT}QJwjBJ'\*Z'IUK_lQ]@'=
    R975x@l<;OWTEZ7nK_2re2,~_jPOtMWXTG~ToEjVmC$J=;m'1DrxG]AH}{p[<#YiIXs2spE=ax=D
    K_RoA*DPgmVU5HoJm<YIk=CwZ5>\!F5i3p]D>X$eG1nOT*|em7~2RTZdI<VIw{^BP1iH<6+H^ejR
    RI3Gs<']^e1<UTn7xTru[pY\wrrHBC+U8=5WG5\Cn1AQ+ziA;_,YWe;[uQ~+1n*x]3e7QMo},Tap
    7u^VpuS',,CxxmB5~V3tXp5}R@]jcI,'_,#Bu-T{,[wneB{+<lmEpE~5]?[5Os[?Qc'Xa?r57X{A
    W^^DOTKORGUsH+)erB.xB&FZU3Aoe>KI+J^la[G6e-]7wwU@#arl_o[@?5=GvE\]?]G'eHB}jvJD
    x=v-)gm7RJ|Yru1iUY}aQKD!j{Ab2E>xs)[WAC&oMIXQa<_n;iwmmEKoB5Tx_euj\-=Yu-Ni5?=_
    T~5^>r*Z$2,kw2R:,s{K\Q<j]oI^O[vk>zOEv\xCK'B*^~r}Y;CEDD>\CCQ~rwO]l=@rUrT+*r^r
    #QQ]_rwYBwl1q\mFeTIW<{QmO?Y\OHYI[;Hr#]IT7VXE$rAr%?t)!hUER=>7T;R_s[lkjwGXpY*i
`endprotected
//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin
`protected

    MTI!#]WVIWUKku*O'{YwOo7=@\7^]<wJBy?Yt[:~]"!HIueQ'#-x;uUz(Q;2KuYCI|=I-J[XWkM-
    {AC@X=pgaap<+1$'Q,AmOoXA31,['>Kj^-1V-]-]_ipHj'As1+B>w[[sB;&}ZEW]G$w{,ACH5~[z
    mvsDK_-NF.GmunCJ-WWo_,2CYH,e>*<QE-~1A-R<o*iGupgpIU?<C=m]GJHUXZGsXUo*Ciza=B?2
    5-_~l#&%@<-1W1<zF\$pu,<Y#Hv<BEU{aHn~Zm\vW]$U?[75Yq5rC_'#A#DxzDPo*~jHR<GHBjwZ
    o~[*#IsU>Yua'ACI+>sx@x;}]Tm?<Bn'3Z!K]wwuqOkUJ:{R@roQ3p\z,@CR{HlBC?<II[>GZxEa
    {HRxsBa7s~AD+]XsBu/-NN$@BHZ=raKn<kI!KjrA1OpsOw?e]j+\?_GIB^XjQ[F{*<xC":1Wxa~5
    @*2+@!i,#Z&1I2kppGksQoi@$p-zz}+Vn2!XG0TexrHAxuT[QrFK[D@TaHuEx#Q$W@oxB<37Eok^
    }ikZ1{zIR#[]W<77ZUBH=oxO<z3C}$^xG#wpW,IG_?;;ET#AO8I5RnJYBrV'G$_d;s+#<'WQ,~rs
    u7rm1Vs]B7Q7B>rAe7X~C/R^JlX]YJ,_~-BV*IUQuUfHC8.Pjzw}(Tr[T}W25p/Y\#pM%4v3K_X,
    C;EemBx~DmYaEw;'CTTT7T[{r?uVls]@;$SZ,{CWz;~-,>!^;veK}KG(5$uO'XY]CC^I^vvlX^1$
    r';Z'&;BeCU*$K<Y+Go-eEKrXpb1TrQG<J^SJDiK_AuCIYjm\H{'i7llREVm#{W3wYTZ2,X!FQQ^
    ^q&$?n?8$KTBB3~?,^,vxB'R$*@7<ET^~^GuZYU}FH<Tp~rsY$;2$K|=HQG[Ee{Kx,py>>xa2T{3
    pm_nRUOpQBawaY\[~lZ?em,=^UlzH{UE=sXjT};-rl=\H_35}TOBBzjBpW'#K]K;QB@eKC,?Z5wv
    HaueR9({{DCUx[Jw]D;Q<oun1<uZT^nl7kv?vw,7AH3_joD+Ym$$[u>djTV~,CO[y;$vTe<Az(AU
    @Ja{QBC{-j^UlTuRp!72],W-HHvxrB3V^@52TGpeVGk5r\us[]H+]$9j=R,D@^#njkB~VzljQJB=
    B$5/=>oWjU8'B[E*]eJ^E#ailwEIxuJ0o>=}zQju{w+*oEzI4E<G_ra*pr*]mnYw?;<aZ[Dc^v{~
    <wo<wxV$yvZ_#BI=$Y+O3p!{[ZI3+nz*iu<s\vsOx\\lCie!jQxaaGTwBl<ru&gvICT]X]iOa!'V
    w]i'R{$[>Om,@Xu*pIR7B175jrs/|_j>Q_To}D*zO\$'HFu{{XsAG5H\3Tocb;zo#T>~-%x'a^Uj
    Z]J'+I]e+,j)pzXC}zuuB7W{LzjXugER{!*x!m:j,C#[UTO7?emJ<-{e]+2oU;TnYOa_1+kPO-!}
    1*K{]^e1wXKZjY]'ssjp#O<~Qv1KU[J}Z-ZJuUVlFqDKXO,Z=Ugl=K5sVQlTV?aT7l!l-DElH<eB
    I^$x^Ar]zeR<O+[n}7sXp[BlX~,^pvkT$IAr-YusHEl'xDO\[oljje@1!=$-D++n$auIlmG{Rw*C
    3=}V*ipH1_OJaz_K7z-sO3Dse<z2w$J:tWhB?uJ\};xzQm]Vi*JmX5@onm<DpG]VIGlm=Am{VK?b
    Os5_}JU<*VD[->}vU[3rcDw>As$~uoeJW]w\x]yw,>1E;IHeo15vGu?5uouYOiV5kY=~n^^~}[xV
    E]K\"G+DE!eY[zj]W1_lJ$w*-^P',5,(r*\_3Hw-LJzpH;r{Tur*]Z>O!OpAo1HG7xDD2']x^Q>^
    x{5}5"k>sjQ}pQfzXmj2Ujx,jW}'[*YIkJk2O?,2[~/v~o+)sloO,i-~o[,aie,G1=>HpR~D]1,'
    B_!>XLC+Rs*{3;TC-R4u7Q#j@p!zX(OTm[sT~Ba}zk1$!-Hp_oGVw26ezezeIoQ8}uK*VZAD3YI3
    u=xU:-,nXfh#[3r],~zQKI^s[OOv4o]B+2o'j[l_$yP,_21<jiQ1Y?7Y^lI_jJE?o}RH73Y6_\?\
    BATX!1uvr1Up"$E<Z:5H{k[TGT-IaTC72xV{1Vvi_QKaZvrY}$QOrT<<RaciYUs[m;QZX{!KUqBp
    _~#a>l\jH;{]r![jmUslj<jrQ!;$}+7}[X|+z~HrBjev1,Z25,krJ2\7_jI}=OHZDCjIA<soiRB*
    >=j^UriIZAY+-QRjJ\UjA~AzuR_{=UE^zG*lUY,5jVl?A{nPl@Ds<Ca,?eZzH<2wQkG1r}3[*JeQ
    K}12r^\?BC<$7up@jWO>Eq1k_n;{ToomD@}u>[-r[@E+ZQ;G~Z#XrDvxV}su,,f[A'mu>vs)Zox,
    fErJ'lpCKER'CU}[A6[@]]>D#'luC\Ouoj9V]r7Ii2;55-Ys#*Tp>z~;=B3=WRvn$U@Vo<[Xwzoc
    JD'E7arY-$$?BIj#7xxRKU~_]3Up$msn}OJl]}I,R'Dsk__plX+G"4Da1i!R~G{+w#e#PrDEZ]ma
    rlur5uCB$IAn_5+A7{wX_R^m-$=mp,e,jT'VaB]7UTO#^)nDz~1A2-j~KV+I^5M:\*>{ut}r?_y2
    rjaW,{u}<TQ*3r^e[xl^kT'Y@QI+DJ@{z7j=iwe#\o~-z,I6Tv1~C_w}q;aeDe;uQmR-^p_Zw!E[
    mB#EKzT!;$$A[2G_v!rkl3YRH#oT]gRoK[$f}*!\k+\@nVKK["@>vnx_ZR
`endprotected
//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin
`protected

    MTI!#-<Y-}pA><Bx2_v'5u-ZxX7m'zr\~j_eW=;7z=s"[B?W,l_uVxW];VV[1mCku[CC:a7-$^12
    wm$C]v--s~{BBY6+1$'Q,AmOoXA31,['>Kj^-1V-]H]H<C;jxmzeD^mmp~@VnjK'IK+]?$I&AUZ[
    p$k1XAY^RW;5znBRNK}oRvERGRRs<kAG~n'vJAET=5KwaO5;K5p[7QwJ#EH1O6HUV~j\5lDel31B
    {}KY_Kd?ORKb:J5,A7pROGBr?isnpzA*\!xB[g3<D7i'C{-YI3_9]kHbBlVT!XRTAOmj#]^]'4B}
    ^ZK[|7?{J=;EjZ{DJ\A_w_Wjz!X^~*2<RHs[i[+JRz-B]~7~e[eBC|G^Yl'urm_H'$3=#x>5<g7V
    }@t3]k@'GW+2ED3JseR=W+[z;O;p\[W_1m',v-=<H\B#YW>nwJ{W[_s!>2e]TT-V{o\C\,!B>Wn1
    RpH!D9aY~^,Ei$EwQ!xI*'R$R#Q'Az^Q>Zw{Yzdu*$r2vD3^?Ck1,7Y?]+jbK[*DAsGK/7!uYIp[
    *HTe!6BT3slaEJ>x983V>]d@R~BJ+Ks$I,x>=@a5DD]YKo1FoiA>uD71;Ynm$-=itFX=^sUr'
`endprotected
//pragma protect end
//pragma protect
//pragma protect begin
`protected

    MTI!#vk7#*[E[IH*xr?WDXoVD}U]u}'%5!-5Fqg~EkTF,T[D>[2\U,?#7\!w=JBvkx-n=-ATUopm
    AXOu<|OZz%lwJ#*+[[o_n=['CW!Ul$HUlIH-BAIz#^^BU7['B>>=i=[?{}XYeBFBFz,!H!YlTf<n
    w[vG3_k<{>&!n5W'BVuj3j$ee><ep,@G{H;\j#[Epx'!'?wxDj~l?z-5K^jFj>QoICkmoTVES>$;
    vrK\?}GOraDQ,nj<p+YG][j}nu]*Rhl|Q\G]LD~Iis5?x@sEE_E{=O'uzJ7#G~=I'_jil~'HE7*w
    *[@]<]T$*e*Q_}^ROKw3vm$i#~x<ZoVZA\QTw'{wJ'2Bp~zZU$?DRjW7x*OCps==R~R?nV5QDRv1
    r2t$\->B\l2}-pZNY#A?oJGQJH!Ia}*Bns}="3esl,3ARJD?5TT7s{<=ju[uEZ7u#i^O#<,JIk5#
    -?r}2kHuXB,nUt?T,iCiV+3A}i[;T#-^Ia,{Aw&\T~R77K[HBs@=~-^7z$oxB_!*VROE5G\Ga[RO
    v_!Dj[},+sk=ure>UOvJHIB[J[[w>O,}YpDr<v$'W3VpznBBvA~UlrlAz+;Us<,ZA3*rlokE\xZ{
    B;XVWW'$+WQkQ';>5GjBs3o[;7D*=Dm=[E@jB+rY{*2dGUspzlepBAOZW<~uB:BKn,l1$m3=OB8E
    VC}uV*5~v\n#+'}$MHwv!$IDHXal@qH[ZzbrX'izEYG$Br~o?J^L\@{vywo+J1pRsU<x@>VUp$_@
    @l>O,tQau33+ea+|6{wJU5x@r]~;#u]'[Jo;3eGI~Wr@E[OnOIR\3=1*BqBzzO#TE>>E#WoT2={T
    lE^]A*v7VOkX[JiYD$wE#>xe+}!7w[vY?$$[Q@RB7+!s<Qp^1^x;ZQ2pZ7gI+K1m]WE\;W{JX3]m
    }<xr2E$#Ge[V%/=Q~[G<u]s+U~f1T}Ev^H^v^5$x~'O=p7kwY>UE}B>'{HD<,QaBnZvZV}-IioRr
    C_@js^eK1,a2r{T-T-J$Ysaxnm#{lEuROD#?z'Ron3!@$]{CU[xi'Go\R}eCGrXYG7OwG3H*oaB{
    ,C*=u*Ob>D'@v!!JpQ]ew<w]>r~-KaArs,E-R1=COH@#bK5OQQA~W|"lIux"Iu@DTj>7}epo1Y~3
    i}+srDGZo&Gr>^;]E76Wlx!v!'AxxK-{BxGsbl-_En_#~eT-w\zJ>]Du~G@uu,u>BQI<7x'#^R*Z
    ~V!z_N^kW}=1l$8tICkCcx2'w_T[w3njr@7j$%V[wB5l[$_la+,H5jE~^uvV$u!+3V>7!E^zDG=C
    #<C3o@2z,>1$C^^m,I|l@z,,B~k^>K'H+3!wQrw!Hn,[!'?DK}c5ms1dJ}\WrDD=[an<l#![>5w~
    >nnI;roamz>3a(N+wEQuXv}/*>KW\aLe#Cu1s=k*iBi<'I*@vT{%ensW}TKQ7_Q+?<c'ebW-rG=#
    {sN>$?eC[<e.!n~u<SF,RKo-]5>svQ}#EA^JGCT]*YEo>vzC'WWiw~2t].@1\momK3Y3>B<E_U*p
    ~B3^H~<EXzS}?wl8Y~=E_BE\nO=?ekxwj1'Y,\nT75IG_eW[OH[~oCK1F@IjV}'{u7TsrGuH#v>w
    AX{KZOBYoxn}QaoJKrO[@[u\\sj2}pY5*Tws<Jr_iONQp;GUUJpZa!}sHwpm*f(1QTDRIeR}i$xC
    '*]dH+E>b1%@5xi]*oTQS=A]GC@UAp$JK#{-a1\Q*r-[+sYuY^C,wn*^@?lio}rjWW[1,v*mxBZ+
    \|Ernp~XX~b~sW,;\+BezYXYD--B!Ku3*nBQI]Js13O6>H5C^=WZUzvsFV,V5}2,G^Y$>*k1JHnI
    ^3I{Z^sGA${mKu>>Q:1O7^_w;x$\2QH'?}.IX>Vm=#-)v?Q-*+jKv_HOJ,pR;]_Wmn7BI~aELpRG
    o5EClAHv#JD*{VeH@lpG7Q?OIn_VpAn7\#lTBr-{nJzp2glI$O*j1#>Xe{UBv1jXlUqOaW]HeZp:
    wY7;!Q7;xz#J1iUClm1TlJC25uKTiT7u.~j{^VHU\U*Qn}*$Y,J3~O3@HUvnzW^-CzRvI^x21,+]
    J^7$*An2+E-Vsp~uaC?22V@7Z:(~Uo+[W9XQ,x-^D57szUx_,^!U}!.z-I>I'k{E!}'ZEGT5TC@N
    0'_5}\!R\YpJVn1X^_1OK?Op#!^THqw{J7_,=x?<>u{a$UcYQZO#AmsYW-HpZ,;=U'nC<n]{A_?9
    wT*=CQQ3r\K!R1EZtuBuDYuV\E-$ExCZ@;1!ar?=Dwe'<ZjJ7jOT\3R5C+aY\^>nDHG+<C7ARAXz
    ID_U_J}iB+X5+nv7QHEaIJ\!p^T'aT\2@pKeC=IVs!^ITBZQsl-\,YaxzOHo^TB3G}]?,>_}WUzO
    $E*7@uauY@Dr?x;^3*rBGsI**MoT\YY5B<o?Te-wHVr{TBT*imppTm?AH~L1e+mhaavmLrO!+QI=
    H,,e>@x75q'XTkvKGpK*5T/'1{#OJDz+z+{@=#D~*}X^r*?EarsjSV]p}}cJn_Z><IZB3D,KUDn8
    1vr;5alRQa+QIFr?A!ihn,[!&@7CUBw7#Ae>awzmv_^ZZJoK5Fev=GA}+vzIl,Vt,.W$Our_Bx#7
    DO,l7UB1s^ua7X\llOzJrxgA\k}Ia@x5s_B&$_l}OwVVkE?--XD{zj$xD!I-wHDC3OO2Y7DA#XYs
    ?<^o@G>e;}7QlsQKm<{s!,=UwsW_izD~z57?9pAa[u,\i$>x+'*>DE^+ZXO5uX1{Afa{p?\eH_ND
    ~e>jz7-<};+VnYKp-]]d_r$_.e6!\XsIXRne?3OApirQwY3SZV3W>rDv\u-$nX}j=Ri@RGI*IIn?
    1B{lo}#W'Dp-oC\ExpvY3]]=rJs2pJI^wpTHHACOj}UevXWT^uD$iQ#jJ*Dm#hxae3uR_~a${O{+
    DaialiDG-,$X$jl^{2QEw+J>}^}iRvWwDZGZ}_jp27ko>lY#^A<>5p^~r14+>,]HDJ$#Go3$J1OY
    dYmZl<\!@I*Z_WDBE_^;G37a=\}ZC>X-e+vB}U1;pB>o3$6!'i$PVC7<^1o-J&=~\}T'TW~De+Wa
    $TOlTzeveZaO2Jv1Ikye\JG6-lz;B1oYV[^*vN<EI]s{Y+.#]vHBoJ11=C[e#p[$uG<lkJ^=u3s'
    eBj7]+E%!+UIn5VAv}Y{=D{~Kz@Dr]B7],7J+G=w!nvlZI,i}Qr+!j$#WHU1IRn{m1+eX_{n~+51
    !s=QIDUUXz^plZIJP^HzI+vs~XV5{$5m3R?j$xT\ln5QaG2Hp%EaQEjC1YLaG{D<liuF5Yn]]Ank
    ['}[EsY@^d5;a~]BTaE>>xi\{_&!pAXdj7!*YUE,kp=a77[DRvWl[UBY{<E5I'KVp?\wQ]R{vBJ5
    ^Z_*rW[j=2nU5X<xYCAJHa-so7]o[wzm=SwVW[5_@UYW[5ITD[T&aApa+j'u@DT7RVD5w]j=ru,~
    doZu[mOB[^@m-B8RCuu^^IAJRswAEaDvBBCT]}}u<$77D[D=p#R=JuXanVWFqawn+KEe*kQ-j^JG
    ;$k-mkH],V2Y'[lk327^5K'\Y4xv+@!o@[TY-}R>uY~}+@xV$Ie>Qvie5K?XB;MmI--1G<nRu'OR
    Ek+KrT+>w-rIUw3:ZGR{)ovjrs*kszo'j.TBVT[B<!{l>39FoN#H[^@jCpkv@ez*$3$_GoL>1j}-
    CZ<B+K$&*zTD+XlvK<ZK@$-U>CECFBHnolo>Aj[{oq.vYVAbm,+ZEGX+wA3W8>YkrTne!cVNH+jr
    7W1[;l[mX{'[p2_\@Hvaw7
`endprotected
//pragma protect end
//pragma protect
//pragma protect begin
`protected

    MTI!#O=T*6xw}kKz5}Hp1mYsWK[m-lxOaRle'i=#o[|*yQ$-Zi}W+-Ha#XsJ}}g)FG;p$#^<,}@^
    Gm'li}mBz77?@}aJ35/o_n=['CW!Ul$HUlIH-BAIz#^^BU7B3v?~'#ej\e*5{ek/[;^R7Z*_v3~T
    sla@D3Y@73olz15IV7)Q=OB({O?Ermjw*oBrxuD}z^_+=WD{]5k2Y}OiV!YX]s1w_EZ1M^4h/2RD
    7?Um_;*BWs,km#>e[-$2u*Y7JeRv\7VIB=1J@>T,JK}VOrJ*k_U^Y*ZEjI+CY}F]sK[3{vm\|ZYz
    [i<z]2=|Hz@@pTmrXo~U;sm7~T]~aG+l[*_KvTp_BGi[EkxEJn'p}kYi[#JQ\nriB>ooG@zlRV]@
    k7D}A[{>{szk#]~}=<Qkz{3QVW\WADz]G?CDE>B5eOuz=2[[NwX_,pWxGFzKXV>}Q$Y*V+nw,7o-
    OK7mv->j<}Av{pUwEaDx=,ZE#x'23^^Qae\a*1sBQW]I~]JsVk}2D12se~~al7qBQHu,ZKQ[3QZo
    lK?;>'@AI@j"'WskG<ps,<
`endprotected
//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin
`protected

    MTI!#xsA7lADGW-j?o2sA=RC#EPwUsRO\UO51kTU]Oi0iDoUzuxO{p,$Cnq6Fhprxu~RRiIZn^{]
    nKNxLzGC[EfkQ'Be-e]iXa[zx^QI}VCX$sD72[$N!U'wz,3!-^DU!tK5a=/aok#Na>mIO[T=*;V{
    vKDj^KYV}s#~H}2!mD<\C&t6x5{o#{D1rA)#oDx*w+k[4G+vm6Uj+ee#^Y<X1BY[BuTw*J}is*$#
    OsDve[]\E-i_YTC0s#zZY_eAprKs+jG5%cA9'EK?^zJCOx_=-wx*C]3U:uAz]@Ru?_UB-=;=kgR_
    p}XTlX}RWA2qp_X>HOQ~lXn2_jvxX{ZrBROkHVv!\x?U+SZw{TUwPEcD$HTeCZsG3=x#|RC[@EZE
    zUrV>]Dn+AC}-X_r{kXl[c"(!1[sk]o?uE#^D{D~CZxW}1X7g>rm@2]QJWo{mZD{}Ixr{=3aU=4f
    5}KrXvE!?s+OD$>'r:g\l<lq%},#@jCRxa{no75X[_};x'n2e{r3XJD1*~'jW!z@JY?}}*a[JKeD
    {is#2QCAeRR(25P^2>sreY[eTTZdloi$(nY^wC!'
`endprotected
//pragma protect end
//pragma protect
//pragma protect begin
`protected

    MTI!#aQH_~vX7D3xwj7O}a_OA=Xs5,i2?[ma~73Y,x0V@7i,#m!7,'[W}ZE3zm[o!Zncm<=^C!5V
    5kj\VTm[rZ,%lwJ#*+[[o_n=['CW!Ul$HUlIH-BAIz#^^BU7]Gvw>Ri=[?oKhksu]x~Z5Q-$>ogl
    OaUi{n]k_]C}=5#TV_^F#*#5o+x!aY7p~}g7L;$+2\__[5s\xV>E1\e~jEVE~}RQVOIY5kQ<]e\*
    [wa}[]Xa2*a3X^3sYU,DH=&AYQz=zR{7Bk?|[u7^#eTA[];<uT,pU}i-z\DOPT5#kLh}P<eUTv1W
    >B1\]IIZQO,RG}lK50U,C27{-\oE[iCsTJ[?u[Bm*Rv==CDk}i,>l17k7?*E]7{n|o+e{3_llwD#
    _QW>p+I='f,XOi%Ve^HkjRuBG~<[lm+2T1=?eZ7jHOovv3OTHInYX1w1F},11v#Y2ROm$vZOO:Kr
    z7xH>wrOQvE?mevzs{RvT[pTYs_w+w\YQ!QsDi'@[5joJp6$JpAH=J7jln;eK^J2Y[@Q#7$WX]Gz
    K]o1pwHw-K[^5x,|%@sXDiGB1pEEIMx@\7+7@<)3}kn4\WX2qJ<{?:ys\i5aQ{#'=H]51_E@Os?B
    su_<oa~E!mvnRDEw'B}LdKO{XB]\2OO3!9=BSjA=\{1uUjTl~E2>aHC'#x\UD4;a{*7X',U'p,Fl
    \;WGU@\gQcUAAn-CT;KDn=W]!$2-TZ]XHJDY2Xv^jn=#W#i-'pz0JG<amA5pe~sXoCk<oUn^)9lV
    [\Y=k2@7rpy2[C{-r'pE^!'p+aTKT]prJ=@Q@|Q,xuIH\m'J*XD3IGNEEU#rDE{XY^prMVS8YZn@
    rlR@@aO?=uo?r)I!'^{,K~e_]]novvUE=liV3HV$rao#o{ddEV[,1}IwBxlu7<a!ll,Go_H$qvW$
    $xITEzj!5#alK^un~wXEG\;K;0V*?A[i>u_J1V}%5~$E}K>zZ7J*?-OsOMBA!sX$Z<'>3wn\?@N^
    J${/@njZsj!XYj?EG~$^BeAC7Jvu,!-D'r+]wQjx5777RYvD7XQxx3x,pQVo}[iu9*a*uW_]p(!E
    lp"G_[uwAI]KxXR-I_IDpkOuXIJrA2>A[AzD#oCRa,C$eau[rY'~rH]^X75-xm]}I-sv15eQ;z5E
    zI,'X-szpOB,G$[okDe8oT$'wo$I2GOoo;@?6xJ'Q/kBRuw[DES'1-zaj13W$*$,u1O'?eBUUz-8
    \[l3XrE\jTsoB^-o\),^U}<ox~kAEx,0#Qv^Txk~i7^~kAJXI_CVP|]rBICC]*5Ok'oWlBHw]2[2
    1sUQvul1+2^VBoA}}_cv7$~jBi7,VeOiE,H{_p=AxOUn\so+5';]G?KlrY@nB,j]3I,q{_u-1Gp#
    iGZjsB{u+5IpK-B[TOwurrD@Xo1Uj$zUp$-2&?vj,)m^r7HzJK;$U<Ka}u7jD!_D'e'^#o6B!Q7F
    551pxTI~~Tr\*gv'KT*_3{74YUsEYZZI7G7]^3esa,e*Pl!Uw5y]CIW<Vwa!|'n@3VH!u_m-san~
    K<j=GpAC@dC-U_v[xac*k$'3]~Zk<+ZA_e@UR>K?,Rs;R'!M*35RB}uj!GwWM*;sWiEn~}wuHWD7
    iYij{*Gz-|zGADRQ']e++Tr[kDm_VUH$T1$k_2$?p@CE{E_uOI"1^R@1OE=.T.*?[D|uC-TP%83l
    p?I>~{Ig$B;a2v^>[\akx$+RD*},@eTEA_}e4z;TV*eDXWwUneDRKj%X]\[}2]{rjA]tE_VB[7VJ
    Bxm@W*3rmqTB=G6h!HOYDXs-$_RI@QZ\,xDZ@5}iJ-{KvIjlBevQ1oZ=jVv5OO@^P%y,^vOE^_B#
    I^e,1+\1BAeuR>$kxV;U>Rjr+s#r\'o!lnTKX$WnUQ3ppxkCvjp0wOY=#e1<B~A--'1?\HY~Y'wz
    3Tu^;H-\<QRV$DA~@o2\,Q12@G\$OAlme-2p^=Is[<w-7!_vEsX;-,,36vj\T5oj~OG6KpV3$[>\
    sUO#Sgx$AuE'aG=&-<Q1po>x'*wvxuVEBX]mU_5Vw=Tm,EnE/AV[-ZQZW,lr],@'Db\,s*tCUQYZ
    x>Oz!CK!Q+!:\B#ZI>Ou;Yzs4Vom}bVeaevs_XY7X^NjX5*hxD*!'aoC^u@U,'TsQ?'~}'o!oQj>
    smR^ZpJ?TGo*VkZ['Aj>5EHptR2-\<\A3'mU@>*}\8TRilxTW+e@D=iSh;C~>T]Za'RH=72Brre+
    ~'O=
`endprotected
//pragma protect end
//pragma protect
//pragma protect begin
`protected

    MTI!#J={>rG;spsO5'e*r,Cn5U+;n,,k7xeUw=3l,e0"^f+sx+*;>Q"EjR[}?,Q2rW@z7;}k5B?~
    [B?I2TX>YT}aap<+1$'Q,AmOoXA31,['>Kj^-1V-]H]H<C;j'AIrZumw<2u*Z1[$mE+]?jI5u$#R
    Z@@GB*#}nuK:u\]pG=wA,l^[{G\*wasXsAf{nrD@E<Zj-I^Js3aE?RuIiUZxK7z:HTE#k6i+sXz$
    w\*32vJGaB@sAEF=_]5k<w~EaZumVYpR~-eT}DT[Cxklx$ik],U(>1oGZe?5!<1r8EQ~!7l}T$ue
    ]h$~[zeJoClvnx)~O!{IUAuTAwGVRUzLBmoiKRik0:G<~1]6kHB'..vH$p(@-E]O<=}[JT2BE3mh
    '!*B$Gr237GpaN$7@k[k1+}'JJ{BTYjAn?Qz*^H]5eb|WzvT,-\m'Q?nD?$v}ZJWHB*Br/G#+}N'
    lZzi5ACzvnrO$=l-wmWgB!$<P"Ba[{',XCKvoQJjC\KExp7,ZUpZ@U}F-\v'fismh353px!j{aA-
    !Y<[YmEHnt>T^=^uOO31+nDEGC)lpvi}.'EROYzujesYmVnlYFoQ~RI2*-OmEAr?Iur\Di#<_oD7
    !Qn5l\^MH-XBcw\X<X{C?6Y}k@pvDZz@m^VQv\IRD$Fy\;X{io5G6|%q]Y1_hgkjD7aeQsW*!2*R
    2[~=C<$!ZEG][#,Qj2'Rv-L}j5=z^Goin!1e7Z;kEE]:BZ{WLg]EKnQo1+r**r%^V1z$E=ai[B[w
    DZV$Ip>{vj[;$z*#G^=7nB_uNrzJB2Y\]vwAQz*1z?GlBzQj*K[w?W*2VR*<mA5^VIDVjX-jr]QG
    *CIllssOJxEO[E<!r~UwIU+Va.iRAj_QAVDI}ZRGoe?D[=Q>ATv[OR!Gr?5rDz$7jJb.>X'!#zw[
    3{Ap_$OiY#E<eB2;Y1m,QYG,IsxAuU][7ekXmIxIo>=$K{ABrvJ?Tr'aCgre,1oC2a\=x~k+YuZY
    ]}1-jX=v5u>$*3lW~aWUA\2[Z\Tsm-k+DRp?v!m_+5TEs!mTOD7@1uh1-<k{j=[e,]ADJeV3I!EV
    WTT$l~QY-{kmtuDuWaEiB'oD[4DxIj27zO'3=k@\D_3z,lz+j1eH;Q7+]B+8G+5{H]#<BpawjzzH
    Hl1#y5TD[R#am=Aoz*&pvDTfizaEKtQDI[X=B;D}u<}v1v[*$J!C$!@snC'^}1IljB&#'X[@=wj=
    ?IuwQAY_nWvDzKuo@,mjBKHKr{oc7$\@uCDYijA=zU2Ino?\R,$xox5QX\C?swW>VDx{>Ul>axE~
    Z-e@DOp?4'ejnE5QlR]UE!UW@]aKE'oskSC7J!DCm7R^O'aAWuviQU-xGjiTVD4>_o3oDX^e7X]e
    e#VA8oXW]C$^#KrVZ'-lW^UeXiEXkKUR~Rp;BDK*VHVv!ON7r-OH]pEZDu#gqn-+~OZH,jGY*[HQ
    }[iDepxz\!>VC{UZzj+>=C[7!}m1j"7u$rO{;W/'5~V[v$pN,[>51n-}H1C!^ko_xK5u?\jpO<lk
    E#BZws<XMpXoTk=epNO*;XzPjsj2-=mGTrow#wQBV?prYv-,I,Aa.I=voUXo{[!6d<<{#~ax;aU_
    _?VW@}TJoInx3*A'Ge'D?Y]vDI2,mWp?YxX5*Gk,UQ5*,IXX',-{Gh"!CG2QeC@'<TW^}DGpi11B
    -l@)EB]D7<R{Wxw\F_rBjB@3Q:uY=]k>E(!w<HviZv!E}i/>wB7QRU+fevo*7~ErEY#p5X\uj'~u
    @puOc;G#;eYWD9.7fp~;}rsGK_arTm]QwKEr>*=1lhgg=Ou_#AQxm1KT%<l5*n^X+o~ArU11#*nI
    ,p{V]l}5BYHVK,UYakaa=[[p1&eloYs}zaZCik~5l+&#TUpvDGm'IDpZQ>Zx!'m1TBG2H~E"'@]O
    vXX>U,r\-}?=piDZo1uDWU'+/J}omwTn=Jnv]C2Jm5VrGu6>{BVOm1V|rEuRzzC,k}1Il?[l5Ok_
    T1@C~CA,]]*Tv5U[I;z2~ln~eKB\lAoG?rC_VcGu7=mY]3[bnH'+{R~RRx@v3zK4wzAeA]^TW^~a
    >X2$WB*mCnQeD<1oo53n^xYVp{,K-j\lxWwTIu6vUxms~[Ym\w}pamHl,B{w,=!3RYDG>raE?[Jv
    RpXQE7#[w[K-w$\WB+Ru[?sSBZ~3GZpY&s5DlHUYWYT@?paQIa<3!:^2*<^HBC[WADz[$IdD>_!+
    ]$rEWVjKtjV*Z<[\x;}u'i]{}]e{7I$p#)&_ZYsmB?[v=;\pzx<5+*;vI-I,r#A<l,_,!;7\~Z=B
    'kCoa@eHxJmGXau!*sKOC>Zj=;o+XjZw7l7k}1rusOuIE7o^-rXICl{5Zo,kX1'xW~;IE<T=Tp=k
    lY}wQm_IKp#vDG}V+OW$]}<zZXKN5Ha;,ajix$],DU5D7,,2AYax^u5UBi5=YY!}^uC=-swoVRw<
    vD]~dGUW@yK\3_->O=<}{-i-^;!]_<ArAQoj-Xw{ACC{;@Vu!Or,Z;_=X=EY73d;r;2*Y1uB37}X
    DUDrDoe[I#JVE?C[!*HIx5C@-_QUeK<G~RE^kxl;OJsB%Yso7?AomlBs;3Ika--OI[<!ujRCs&DY
    B;v<AY~vA~w=np{<T>7[[X_a5]CR?I^!!2E5C$2^?2Y!x,'4%BX]jXT5@kX'XKC'Z^o*^4zU<a=s
    ETC!X^U]=ZlYie7pI+7r5@seQXClRZR@3G)p*To\]^[QH'<[r?{TU]~EQ$J=m'w/-tkY?{ccdx+@
    R_JXGc_\5DAU@rs2Dz*uRm/iLE+-upTWksDH7mY@=]ZvpzUXuD?+se<-7d*?au&W*-U<GJE^2Ga*
    ij*DU{oU<KZ1IxJm\$Uf^3^1#X$@kCsl1B>>Nv*ARKTUeg]uKTCX5=<$T#Xx}I{GGkp@OQu}IYCX
    ]XEYw*U\^}}T;W$2B+@vJ]mGHk#1A<Fz^[lCBI^a,{}r]3}=+N/ID_JLB_ok9K=,YYaaG7V=OzoT
    2=1s^"six@YkX)I2+'6mw_J{G=!<jHG^Ua~J}p[l=>KCzrKjTG-DiBW>Y<ewIU#$3eoJsJR@vmwi
    Dl,D,rlxB@B_wwY$O}-ap#~${,po[,*m'Tk7VE~]]<Zs2<snjx<*XoT-OuG~Ri=6r*1Z_BWQvXR~
    @ExpX'U7GsBUDz[CjUoXVV+JEJ~HWORZnYA<T1Zjwee@p5Yp}dQ\A?ST>+v@,l30mGX[C,@YCJoO
    a-VZx4oa5;$=]}<w\~HR#RC@!IyYwGV^l$$X^Y=GKm,mvon~\<G'vi1th=?U?[vp;^3-ep!1z?_~
    r$;Hn@D^GvUvBUExKE[K!1m\n'Zo#}'zx_EG;nn3UAT$oOgDl-;$^s>ZXCaWHrUD1+H}#@*7)=!K
    ,D#r>Iok$}RsneC=,
`endprotected
//pragma protect end
