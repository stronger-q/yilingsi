

/**   这里是滑动窗口生成模��?  **/

module BRIEF_WINDOW31_31_1 (
    input                                  i_clk,

    interface_image.i_image                i_image,     //图像输入
    interface_windows.o_window        o_window       //截取滑动窗口后输��?
    );

parameter Pra_Value_Width=8;    //像素深度
localparam Pra_Window_Size=31;  //滑动窗口尺寸

logic               Image_VS_Rising;    //用高电平标记垂直同步上升沿，表示图像帧的��?��?
logic               Image_VS_Falling;   //用高电平标记垂直同步下降沿，表示图像帧结��?
logic               Image_HS_Rising;    //水平同步上升沿同上，表示��?行图像开��?
logic               Image_HS_Falling;   //水平同步下降��?

logic [15:0]          Counter_Image_VS;
logic [15:0]          Counter_Image_HS;

DVP_Counter u_DVP_Counter (     //加载垂直同步计数器，记录图像处理情况
    .i_clk                   ( i_clk             ),
    .i_dvp_vs                ( i_image.image_vs  ),
    .i_dvp_hs                ( i_image.image_hs  ),

    .o_vs_start              ( Image_VS_Rising   ),
    .o_vs_end                ( Image_VS_Falling  ),
    .o_hs_start              ( Image_HS_Rising   ),
    .o_hs_end                ( Image_HS_Falling  ),
    .o_counter_vs            ( Counter_Image_VS  ),
    .o_counter_hs            ( Counter_Image_HS  )
);

logic [Pra_Window_Size-2:0]            FIFO_Full;
logic [Pra_Window_Size-2:0]            FIFO_Empty;
logic [Pra_Window_Size-2:0]            FIFO_WR_Busy;
logic [Pra_Window_Size-2:0]            FIFO_RD_Busy;//efinity doesnt have
logic [10:0]                           FIFO_Read_Count[Pra_Window_Size-2:0];
logic [10:0]                           FIFO_Write_Count[Pra_Window_Size-2:0];
logic [Pra_Window_Size-2:0]            FIFO_Write_En;
logic [Pra_Value_Width-1:0]            FIFO_Write_Data[Pra_Window_Size-2:0];
logic [Pra_Window_Size-2:0]            FIFO_Read_En;
logic [Pra_Value_Width-1:0]            FIFO_Read_Data[Pra_Window_Size-2:0];     //从FIFO中读出来的一行数��?

logic [Pra_Window_Size-1:0]            Flag_Line_Ready;


assign FIFO_Write_En[0]=i_image.image_hs;       //水平同步为高电平时使能FIFO写入
assign FIFO_Write_Data[0]=i_image.image_data;   //为FIFO输入配置像素数据
assign Flag_Line_Ready[0]=1;            //第一行的写入准备标志常设高电��?

logic FIFO_Reset=0;     //复位信号设为低电��?


generate    //生成FIFO_Block块，将图像信号写入和读出FIFO
genvar i;
for (i = 0; i<Pra_Window_Size-1; i++) begin : FIFO_Block       

        FIFO_8_2048_FWFT FIFO_8_2048_FWFT_Line_Buffer_31 (
//EFINITY_TEST
//        .a_rst_i(FIFO_Reset),                     
//        .wr_clk_i(i_clk),                
//        .rd_clk_i(i_clk),                

//        .wr_en_i(FIFO_Write_En[i]),                  
//        .wdata(FIFO_Write_Data[i]),                     
//        .rd_en_i(FIFO_Read_En[i]),                
//        .rdata(FIFO_Read_Data[i]),                    

//        .full_o(FIFO_Full[i]),                    
//        .empty_o(FIFO_Empty[i]),                  
//        .rd_datacount_o(FIFO_Read_Count[i]),  
//        .wr_datacount_o(FIFO_Write_Count[i]),  
//        .rst_busy(FIFO_WR_Busy[i])

//VIVADO_TEST
        .a_rst_i(FIFO_Reset),            // input wire rst
        .wr_clk_i(i_clk),                // input wire wr_clk
        .rd_clk_i(i_clk),                // input wire rd_clk

        .wr_en_i(FIFO_Write_En[i]),                  // input wire wr_en
        .wdata(FIFO_Write_Data[i]),                      // input wire [7 : 0] din
        .rd_en_i(FIFO_Read_En[i]),                  // input wire rd_en
        .rdata(FIFO_Read_Data[i]),                    // output wire [7 : 0] dout

        .full_o(FIFO_Full[i]),                    // output wire full
        .empty_o(FIFO_Empty[i]),                  // output wire empty
        .rd_datacount_o(FIFO_Read_Count[i]),  // output wire [10 : 0] rd_data_count
        .wr_datacount_o(FIFO_Write_Count[i])  // output wire [10 : 0] wr_data_count
        );
   

assign FIFO_Read_En[i]=Flag_Line_Ready[i+1]&i_image.image_hs;       //i+1行数据准备好，并且当前行��?始时，允许从FIFIO中读取数��?

end
endgenerate

generate
genvar j;
for (j = 1; j<Pra_Window_Size-1; j++) begin : Always_Blaock

always @(posedge i_clk)
begin
    if(Image_VS_Rising)     
    begin
        Flag_Line_Ready[j]<=0;      //出现垂直同步信号上升沿时，原先的写入准备标志置零
    end
    else if(Image_HS_Falling==1'b1 && FIFO_Read_Count[j-1]>0)   //else，前��?行的水平同步下降沿出现，和FIFO读取计数不为零，即数据读取完成时
    begin
        Flag_Line_Ready[j]<=1;      //此时将下��?行的写入准备标志设为高电平，即允许读取数��?
    end
    else
    begin
        Flag_Line_Ready[j]<=Flag_Line_Ready[j];     //否则下一行的写入准备标志不变
    end
end


if(Pra_Window_Size==2) begin
    //空的
end
else begin
    assign FIFO_Write_En[j]=FIFO_Read_En[j-1];
    assign FIFO_Write_Data[j]=FIFO_Read_Data[j-1];      //将数据从第j-1行搬运到第j��?
end


end
endgenerate


//为滑动窗口数据准备寄存器
//每个数组储存��?列的像素数据，每个数组元素代表一个像��?
logic [Pra_Value_Width-1:0]        Window_Data_00_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_01_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_02_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_03_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_04_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_05_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_06_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_07_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_08_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_09_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_10_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_11_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_12_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_13_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_14_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_15_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_16_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_17_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_18_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_19_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_20_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_21_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_22_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_23_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_24_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_25_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_26_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_27_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_28_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_29_XX[Pra_Window_Size-1:0];
logic [Pra_Value_Width-1:0]        Window_Data_30_XX[Pra_Window_Size-1:0];



generate        //生成Window_Block块，将每��?行的数据移动到下��?行，实现窗口滑动
genvar k;
for (k = 0; k<Pra_Window_Size-1; k++) begin : Window_Block
    always @(posedge i_clk)
    begin
        Window_Data_00_XX[k+1]<=Window_Data_00_XX[k];
        Window_Data_01_XX[k+1]<=Window_Data_01_XX[k];
        Window_Data_02_XX[k+1]<=Window_Data_02_XX[k];
        Window_Data_03_XX[k+1]<=Window_Data_03_XX[k];
        Window_Data_04_XX[k+1]<=Window_Data_04_XX[k];
        Window_Data_05_XX[k+1]<=Window_Data_05_XX[k];
        Window_Data_06_XX[k+1]<=Window_Data_06_XX[k];
        Window_Data_07_XX[k+1]<=Window_Data_07_XX[k];
        Window_Data_08_XX[k+1]<=Window_Data_08_XX[k];
        Window_Data_09_XX[k+1]<=Window_Data_09_XX[k];
        Window_Data_10_XX[k+1]<=Window_Data_10_XX[k];
        Window_Data_11_XX[k+1]<=Window_Data_11_XX[k];
        Window_Data_12_XX[k+1]<=Window_Data_12_XX[k];
        Window_Data_13_XX[k+1]<=Window_Data_13_XX[k];
        Window_Data_14_XX[k+1]<=Window_Data_14_XX[k];
        Window_Data_15_XX[k+1]<=Window_Data_15_XX[k];
        Window_Data_16_XX[k+1]<=Window_Data_16_XX[k];
        Window_Data_17_XX[k+1]<=Window_Data_17_XX[k];
        Window_Data_18_XX[k+1]<=Window_Data_18_XX[k];
        Window_Data_19_XX[k+1]<=Window_Data_19_XX[k];
        Window_Data_20_XX[k+1]<=Window_Data_20_XX[k];
        Window_Data_21_XX[k+1]<=Window_Data_21_XX[k];
        Window_Data_22_XX[k+1]<=Window_Data_22_XX[k];
        Window_Data_23_XX[k+1]<=Window_Data_23_XX[k];
        Window_Data_24_XX[k+1]<=Window_Data_24_XX[k];
        Window_Data_25_XX[k+1]<=Window_Data_25_XX[k];
        Window_Data_26_XX[k+1]<=Window_Data_26_XX[k];
        Window_Data_27_XX[k+1]<=Window_Data_27_XX[k];
        Window_Data_28_XX[k+1]<=Window_Data_28_XX[k];
        Window_Data_29_XX[k+1]<=Window_Data_29_XX[k];
        Window_Data_30_XX[k+1]<=Window_Data_30_XX[k];
    end
end

endgenerate


//将FIFO中读取出的最新一行数据赋值给滑动窗口的第��?行，实现数据更新
assign Window_Data_00_XX[0]=FIFO_Read_Data[Pra_Window_Size-2];
assign Window_Data_01_XX[0]=FIFO_Read_Data[Pra_Window_Size-3];
assign Window_Data_02_XX[0]=FIFO_Read_Data[Pra_Window_Size-4];
assign Window_Data_03_XX[0]=FIFO_Read_Data[Pra_Window_Size-5];
assign Window_Data_04_XX[0]=FIFO_Read_Data[Pra_Window_Size-6];
assign Window_Data_05_XX[0]=FIFO_Read_Data[Pra_Window_Size-7];
assign Window_Data_06_XX[0]=FIFO_Read_Data[Pra_Window_Size-8];
assign Window_Data_07_XX[0]=FIFO_Read_Data[Pra_Window_Size-9];
assign Window_Data_08_XX[0]=FIFO_Read_Data[Pra_Window_Size-10];
assign Window_Data_09_XX[0]=FIFO_Read_Data[Pra_Window_Size-11];
assign Window_Data_10_XX[0]=FIFO_Read_Data[Pra_Window_Size-12];
assign Window_Data_11_XX[0]=FIFO_Read_Data[Pra_Window_Size-13];
assign Window_Data_12_XX[0]=FIFO_Read_Data[Pra_Window_Size-14];
assign Window_Data_13_XX[0]=FIFO_Read_Data[Pra_Window_Size-15];
assign Window_Data_14_XX[0]=FIFO_Read_Data[Pra_Window_Size-16];
assign Window_Data_15_XX[0]=FIFO_Read_Data[Pra_Window_Size-17];
assign Window_Data_16_XX[0]=FIFO_Read_Data[Pra_Window_Size-18];
assign Window_Data_17_XX[0]=FIFO_Read_Data[Pra_Window_Size-19];
assign Window_Data_18_XX[0]=FIFO_Read_Data[Pra_Window_Size-20];
assign Window_Data_19_XX[0]=FIFO_Read_Data[Pra_Window_Size-21];
assign Window_Data_20_XX[0]=FIFO_Read_Data[Pra_Window_Size-22];
assign Window_Data_21_XX[0]=FIFO_Read_Data[Pra_Window_Size-23];
assign Window_Data_22_XX[0]=FIFO_Read_Data[Pra_Window_Size-24];
assign Window_Data_23_XX[0]=FIFO_Read_Data[Pra_Window_Size-25];
assign Window_Data_24_XX[0]=FIFO_Read_Data[Pra_Window_Size-26];
assign Window_Data_25_XX[0]=FIFO_Read_Data[Pra_Window_Size-27];
assign Window_Data_26_XX[0]=FIFO_Read_Data[Pra_Window_Size-28];
assign Window_Data_27_XX[0]=FIFO_Read_Data[Pra_Window_Size-29];
assign Window_Data_28_XX[0]=FIFO_Read_Data[Pra_Window_Size-30];
assign Window_Data_29_XX[0]=FIFO_Read_Data[Pra_Window_Size-31];
assign Window_Data_30_XX[0]=i_image.image_data;


logic Flag_Pixel_Ready;

always @(posedge i_clk)
begin
    if(Image_VS_Rising)
    begin
        Flag_Pixel_Ready<=0;        //当新的图像帧��?始时，像素准备标志置0
    end
    else if(Counter_Image_HS>=Pra_Window_Size-2)
    begin
        Flag_Pixel_Ready<=1;        //水平同步计数值到��?29，即该图像帧处理完成时，像素准备标志��?1
    end
    else
    begin
        Flag_Pixel_Ready<=0;
    end
end

assign o_window.image_vs=i_image.image_vs;      //
assign o_window.image_hs=i_image.image_hs;      //这两行接驳垂直与水平同步信号至输��?
assign o_window.image_en=i_image.image_hs&Flag_Line_Ready[Pra_Window_Size-1]&Flag_Pixel_Ready;
    //��?有准备标志都��?1时，允许图像输出


    //以下代码将每个滑动窗口像素数据接驳至输出端口
assign
 o_window.window_00[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_00[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_01[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_02[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_03[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_04[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_05[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_06[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_07[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_08[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_09[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_10[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_11[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_12[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_13[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_14[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_15[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_16[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_17[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_18[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_19[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_20[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_21[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_22[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_23[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_24[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_25[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_26[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_27[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_28[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_29[30] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[00] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[01] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[02] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[03] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[04] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[05] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[06] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[07] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[08] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[09] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[10] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[11] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[12] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[13] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[14] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[15] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[16] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[17] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[18] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[19] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[20] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[21] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[22] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[23] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[24] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[25] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[26] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[27] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[28] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[29] = Window_Data_00_XX[Pra_Window_Size-1];
assign
 o_window.window_30[30] = Window_Data_00_XX[Pra_Window_Size-1];



endmodule
